`timescale 1 ns/100 ps
// Version: v12.5 12.900.10.16


module miv_rv32_ram_singleport_lp_ecc(
       W_DATA,
       R_DATA,
       W_ADDR,
       R_ADDR,
       W_EN,
       R_EN,
       CLK,
       SB_CORRECT,
       DB_DETECT
    );
parameter RAM_DEPTH = 32'h4000;   // Max depth 256KB

input  [31:0] W_DATA;
output [31:0] R_DATA;
input  [15:0] W_ADDR;
input  [15:0] R_ADDR;
input  W_EN;
input  R_EN;
input  CLK;
output SB_CORRECT;
output DB_DETECT;

    wire [31:0] int_R_DATA_TEMPR0  , sel_R_DATA_TEMPR0  ,
                int_R_DATA_TEMPR1  , sel_R_DATA_TEMPR1  ,
                int_R_DATA_TEMPR2  , sel_R_DATA_TEMPR2  ,
                int_R_DATA_TEMPR3  , sel_R_DATA_TEMPR3  ,
                int_R_DATA_TEMPR4  , sel_R_DATA_TEMPR4  ,
                int_R_DATA_TEMPR5  , sel_R_DATA_TEMPR5  ,
                int_R_DATA_TEMPR6  , sel_R_DATA_TEMPR6  ,
                int_R_DATA_TEMPR7  , sel_R_DATA_TEMPR7  ,
                int_R_DATA_TEMPR8  , sel_R_DATA_TEMPR8  ,
                int_R_DATA_TEMPR9  , sel_R_DATA_TEMPR9  ,
                int_R_DATA_TEMPR10 , sel_R_DATA_TEMPR10 ,
                int_R_DATA_TEMPR11 , sel_R_DATA_TEMPR11 ,
                int_R_DATA_TEMPR12 , sel_R_DATA_TEMPR12 ,
                int_R_DATA_TEMPR13 , sel_R_DATA_TEMPR13 ,
                int_R_DATA_TEMPR14 , sel_R_DATA_TEMPR14 ,
                int_R_DATA_TEMPR15 , sel_R_DATA_TEMPR15 ,
                int_R_DATA_TEMPR16 , sel_R_DATA_TEMPR16 ,
                int_R_DATA_TEMPR17 , sel_R_DATA_TEMPR17 ,
                int_R_DATA_TEMPR18 , sel_R_DATA_TEMPR18 ,
                int_R_DATA_TEMPR19 , sel_R_DATA_TEMPR19 ,
                int_R_DATA_TEMPR20 , sel_R_DATA_TEMPR20 ,
                int_R_DATA_TEMPR21 , sel_R_DATA_TEMPR21 ,
                int_R_DATA_TEMPR22 , sel_R_DATA_TEMPR22 ,
                int_R_DATA_TEMPR23 , sel_R_DATA_TEMPR23 ,
                int_R_DATA_TEMPR24 , sel_R_DATA_TEMPR24 ,
                int_R_DATA_TEMPR25 , sel_R_DATA_TEMPR25 ,
                int_R_DATA_TEMPR26 , sel_R_DATA_TEMPR26 ,
                int_R_DATA_TEMPR27 , sel_R_DATA_TEMPR27 ,
                int_R_DATA_TEMPR28 , sel_R_DATA_TEMPR28 ,
                int_R_DATA_TEMPR29 , sel_R_DATA_TEMPR29 ,
                int_R_DATA_TEMPR30 , sel_R_DATA_TEMPR30 ,
                int_R_DATA_TEMPR31 , sel_R_DATA_TEMPR31 ,
                int_R_DATA_TEMPR32 , sel_R_DATA_TEMPR32 ,
                int_R_DATA_TEMPR33 , sel_R_DATA_TEMPR33 ,
                int_R_DATA_TEMPR34 , sel_R_DATA_TEMPR34 ,
                int_R_DATA_TEMPR35 , sel_R_DATA_TEMPR35 ,
                int_R_DATA_TEMPR36 , sel_R_DATA_TEMPR36 ,
                int_R_DATA_TEMPR37 , sel_R_DATA_TEMPR37 ,
                int_R_DATA_TEMPR38 , sel_R_DATA_TEMPR38 ,
                int_R_DATA_TEMPR39 , sel_R_DATA_TEMPR39 ,
                int_R_DATA_TEMPR40 , sel_R_DATA_TEMPR40 ,
                int_R_DATA_TEMPR41 , sel_R_DATA_TEMPR41 ,
                int_R_DATA_TEMPR42 , sel_R_DATA_TEMPR42 ,
                int_R_DATA_TEMPR43 , sel_R_DATA_TEMPR43 ,
                int_R_DATA_TEMPR44 , sel_R_DATA_TEMPR44 ,
                int_R_DATA_TEMPR45 , sel_R_DATA_TEMPR45 ,
                int_R_DATA_TEMPR46 , sel_R_DATA_TEMPR46 ,
                int_R_DATA_TEMPR47 , sel_R_DATA_TEMPR47 ,
                int_R_DATA_TEMPR48 , sel_R_DATA_TEMPR48 ,
                int_R_DATA_TEMPR49 , sel_R_DATA_TEMPR49 ,
                int_R_DATA_TEMPR50 , sel_R_DATA_TEMPR50 ,
                int_R_DATA_TEMPR51 , sel_R_DATA_TEMPR51 ,
                int_R_DATA_TEMPR52 , sel_R_DATA_TEMPR52 ,
                int_R_DATA_TEMPR53 , sel_R_DATA_TEMPR53 ,
                int_R_DATA_TEMPR54 , sel_R_DATA_TEMPR54 ,
                int_R_DATA_TEMPR55 , sel_R_DATA_TEMPR55 ,
                int_R_DATA_TEMPR56 , sel_R_DATA_TEMPR56 ,
                int_R_DATA_TEMPR57 , sel_R_DATA_TEMPR57 ,
                int_R_DATA_TEMPR58 , sel_R_DATA_TEMPR58 ,
                int_R_DATA_TEMPR59 , sel_R_DATA_TEMPR59 ,
                int_R_DATA_TEMPR60 , sel_R_DATA_TEMPR60 ,
                int_R_DATA_TEMPR61 , sel_R_DATA_TEMPR61 ,
                int_R_DATA_TEMPR62 , sel_R_DATA_TEMPR62 ,
                int_R_DATA_TEMPR63 , sel_R_DATA_TEMPR63 ,
                int_R_DATA_TEMPR64 , sel_R_DATA_TEMPR64 ,
                int_R_DATA_TEMPR65 , sel_R_DATA_TEMPR65 ,
                int_R_DATA_TEMPR66 , sel_R_DATA_TEMPR66 ,
                int_R_DATA_TEMPR67 , sel_R_DATA_TEMPR67 ,
                int_R_DATA_TEMPR68 , sel_R_DATA_TEMPR68 ,
                int_R_DATA_TEMPR69 , sel_R_DATA_TEMPR69 ,
                int_R_DATA_TEMPR70 , sel_R_DATA_TEMPR70 ,
                int_R_DATA_TEMPR71 , sel_R_DATA_TEMPR71 ,
                int_R_DATA_TEMPR72 , sel_R_DATA_TEMPR72 ,
                int_R_DATA_TEMPR73 , sel_R_DATA_TEMPR73 ,
                int_R_DATA_TEMPR74 , sel_R_DATA_TEMPR74 ,
                int_R_DATA_TEMPR75 , sel_R_DATA_TEMPR75 ,
                int_R_DATA_TEMPR76 , sel_R_DATA_TEMPR76 ,
                int_R_DATA_TEMPR77 , sel_R_DATA_TEMPR77 ,
                int_R_DATA_TEMPR78 , sel_R_DATA_TEMPR78 ,
                int_R_DATA_TEMPR79 , sel_R_DATA_TEMPR79 ,
                int_R_DATA_TEMPR80 , sel_R_DATA_TEMPR80 ,
                int_R_DATA_TEMPR81 , sel_R_DATA_TEMPR81 ,
                int_R_DATA_TEMPR82 , sel_R_DATA_TEMPR82 ,
                int_R_DATA_TEMPR83 , sel_R_DATA_TEMPR83 ,
                int_R_DATA_TEMPR84 , sel_R_DATA_TEMPR84 ,
                int_R_DATA_TEMPR85 , sel_R_DATA_TEMPR85 ,
                int_R_DATA_TEMPR86 , sel_R_DATA_TEMPR86 ,
                int_R_DATA_TEMPR87 , sel_R_DATA_TEMPR87 ,
                int_R_DATA_TEMPR88 , sel_R_DATA_TEMPR88 ,
                int_R_DATA_TEMPR89 , sel_R_DATA_TEMPR89 ,
                int_R_DATA_TEMPR90 , sel_R_DATA_TEMPR90 ,
                int_R_DATA_TEMPR91 , sel_R_DATA_TEMPR91 ,
                int_R_DATA_TEMPR92 , sel_R_DATA_TEMPR92 ,
                int_R_DATA_TEMPR93 , sel_R_DATA_TEMPR93 ,
                int_R_DATA_TEMPR94 , sel_R_DATA_TEMPR94 ,
                int_R_DATA_TEMPR95 , sel_R_DATA_TEMPR95 ,
                int_R_DATA_TEMPR96 , sel_R_DATA_TEMPR96 ,
                int_R_DATA_TEMPR97 , sel_R_DATA_TEMPR97 ,
                int_R_DATA_TEMPR98 , sel_R_DATA_TEMPR98 ,
                int_R_DATA_TEMPR99 , sel_R_DATA_TEMPR99 ,
                int_R_DATA_TEMPR100, sel_R_DATA_TEMPR100,
                int_R_DATA_TEMPR101, sel_R_DATA_TEMPR101,
                int_R_DATA_TEMPR102, sel_R_DATA_TEMPR102,
                int_R_DATA_TEMPR103, sel_R_DATA_TEMPR103,
                int_R_DATA_TEMPR104, sel_R_DATA_TEMPR104,
                int_R_DATA_TEMPR105, sel_R_DATA_TEMPR105,
                int_R_DATA_TEMPR106, sel_R_DATA_TEMPR106,
                int_R_DATA_TEMPR107, sel_R_DATA_TEMPR107,
                int_R_DATA_TEMPR108, sel_R_DATA_TEMPR108,
                int_R_DATA_TEMPR109, sel_R_DATA_TEMPR109,
                int_R_DATA_TEMPR110, sel_R_DATA_TEMPR110,
                int_R_DATA_TEMPR111, sel_R_DATA_TEMPR111,
                int_R_DATA_TEMPR112, sel_R_DATA_TEMPR112,
                int_R_DATA_TEMPR113, sel_R_DATA_TEMPR113,
                int_R_DATA_TEMPR114, sel_R_DATA_TEMPR114,
                int_R_DATA_TEMPR115, sel_R_DATA_TEMPR115,
                int_R_DATA_TEMPR116, sel_R_DATA_TEMPR116,
                int_R_DATA_TEMPR117, sel_R_DATA_TEMPR117,
                int_R_DATA_TEMPR118, sel_R_DATA_TEMPR118,
                int_R_DATA_TEMPR119, sel_R_DATA_TEMPR119,
                int_R_DATA_TEMPR120, sel_R_DATA_TEMPR120,
                int_R_DATA_TEMPR121, sel_R_DATA_TEMPR121,
                int_R_DATA_TEMPR122, sel_R_DATA_TEMPR122,
                int_R_DATA_TEMPR123, sel_R_DATA_TEMPR123,
                int_R_DATA_TEMPR124, sel_R_DATA_TEMPR124,
                int_R_DATA_TEMPR125, sel_R_DATA_TEMPR125,
                int_R_DATA_TEMPR126, sel_R_DATA_TEMPR126,
                int_R_DATA_TEMPR127, sel_R_DATA_TEMPR127;

    wire [127:0] int_SB_CORRECT_NG, sel_SB_CORRECT_NG,
                 int_DB_DETECT_NG, sel_DB_DETECT_NG,
                 ACCESS_BUSY;
	
    assign sel_R_DATA_TEMPR0   = (RAM_DEPTH > 32'h0   ) ? int_R_DATA_TEMPR0   : 32'b0;
    assign sel_R_DATA_TEMPR1   = (RAM_DEPTH > 32'h200 ) ? int_R_DATA_TEMPR1   : 32'b0;
    assign sel_R_DATA_TEMPR2   = (RAM_DEPTH > 32'h400 ) ? int_R_DATA_TEMPR2   : 32'b0;
    assign sel_R_DATA_TEMPR3   = (RAM_DEPTH > 32'h600 ) ? int_R_DATA_TEMPR3   : 32'b0;
    assign sel_R_DATA_TEMPR4   = (RAM_DEPTH > 32'h800 ) ? int_R_DATA_TEMPR4   : 32'b0;
    assign sel_R_DATA_TEMPR5   = (RAM_DEPTH > 32'hA00 ) ? int_R_DATA_TEMPR5   : 32'b0;
    assign sel_R_DATA_TEMPR6   = (RAM_DEPTH > 32'hC00 ) ? int_R_DATA_TEMPR6   : 32'b0;
    assign sel_R_DATA_TEMPR7   = (RAM_DEPTH > 32'hE00 ) ? int_R_DATA_TEMPR7   : 32'b0;
    assign sel_R_DATA_TEMPR8   = (RAM_DEPTH > 32'h1000) ? int_R_DATA_TEMPR8   : 32'b0;
    assign sel_R_DATA_TEMPR9   = (RAM_DEPTH > 32'h1200) ? int_R_DATA_TEMPR9   : 32'b0;
    assign sel_R_DATA_TEMPR10  = (RAM_DEPTH > 32'h1400) ? int_R_DATA_TEMPR10  : 32'b0;
    assign sel_R_DATA_TEMPR11  = (RAM_DEPTH > 32'h1600) ? int_R_DATA_TEMPR11  : 32'b0;
    assign sel_R_DATA_TEMPR12  = (RAM_DEPTH > 32'h1800) ? int_R_DATA_TEMPR12  : 32'b0;
    assign sel_R_DATA_TEMPR13  = (RAM_DEPTH > 32'h1A00) ? int_R_DATA_TEMPR13  : 32'b0;
    assign sel_R_DATA_TEMPR14  = (RAM_DEPTH > 32'h1C00) ? int_R_DATA_TEMPR14  : 32'b0;
    assign sel_R_DATA_TEMPR15  = (RAM_DEPTH > 32'h1E00) ? int_R_DATA_TEMPR15  : 32'b0;
    assign sel_R_DATA_TEMPR16  = (RAM_DEPTH > 32'h2000) ? int_R_DATA_TEMPR16  : 32'b0;
    assign sel_R_DATA_TEMPR17  = (RAM_DEPTH > 32'h2200) ? int_R_DATA_TEMPR17  : 32'b0;
    assign sel_R_DATA_TEMPR18  = (RAM_DEPTH > 32'h2400) ? int_R_DATA_TEMPR18  : 32'b0;
    assign sel_R_DATA_TEMPR19  = (RAM_DEPTH > 32'h2600) ? int_R_DATA_TEMPR19  : 32'b0;
    assign sel_R_DATA_TEMPR20  = (RAM_DEPTH > 32'h2800) ? int_R_DATA_TEMPR20  : 32'b0;
    assign sel_R_DATA_TEMPR21  = (RAM_DEPTH > 32'h2A00) ? int_R_DATA_TEMPR21  : 32'b0;
    assign sel_R_DATA_TEMPR22  = (RAM_DEPTH > 32'h2C00) ? int_R_DATA_TEMPR22  : 32'b0;
    assign sel_R_DATA_TEMPR23  = (RAM_DEPTH > 32'h2E00) ? int_R_DATA_TEMPR23  : 32'b0;
    assign sel_R_DATA_TEMPR24  = (RAM_DEPTH > 32'h3000) ? int_R_DATA_TEMPR24  : 32'b0;
    assign sel_R_DATA_TEMPR25  = (RAM_DEPTH > 32'h3200) ? int_R_DATA_TEMPR25  : 32'b0;
    assign sel_R_DATA_TEMPR26  = (RAM_DEPTH > 32'h3400) ? int_R_DATA_TEMPR26  : 32'b0;
    assign sel_R_DATA_TEMPR27  = (RAM_DEPTH > 32'h3600) ? int_R_DATA_TEMPR27  : 32'b0;
    assign sel_R_DATA_TEMPR28  = (RAM_DEPTH > 32'h3800) ? int_R_DATA_TEMPR28  : 32'b0;
    assign sel_R_DATA_TEMPR29  = (RAM_DEPTH > 32'h3A00) ? int_R_DATA_TEMPR29  : 32'b0;
    assign sel_R_DATA_TEMPR30  = (RAM_DEPTH > 32'h3C00) ? int_R_DATA_TEMPR30  : 32'b0;
    assign sel_R_DATA_TEMPR31  = (RAM_DEPTH > 32'h3E00) ? int_R_DATA_TEMPR31  : 32'b0;
    assign sel_R_DATA_TEMPR32  = (RAM_DEPTH > 32'h4000) ? int_R_DATA_TEMPR32  : 32'b0;
    assign sel_R_DATA_TEMPR33  = (RAM_DEPTH > 32'h4200) ? int_R_DATA_TEMPR33  : 32'b0;
    assign sel_R_DATA_TEMPR34  = (RAM_DEPTH > 32'h4400) ? int_R_DATA_TEMPR34  : 32'b0;
    assign sel_R_DATA_TEMPR35  = (RAM_DEPTH > 32'h4600) ? int_R_DATA_TEMPR35  : 32'b0;
    assign sel_R_DATA_TEMPR36  = (RAM_DEPTH > 32'h4800) ? int_R_DATA_TEMPR36  : 32'b0;
    assign sel_R_DATA_TEMPR37  = (RAM_DEPTH > 32'h4A00) ? int_R_DATA_TEMPR37  : 32'b0;
    assign sel_R_DATA_TEMPR38  = (RAM_DEPTH > 32'h4C00) ? int_R_DATA_TEMPR38  : 32'b0;
    assign sel_R_DATA_TEMPR39  = (RAM_DEPTH > 32'h4E00) ? int_R_DATA_TEMPR39  : 32'b0;
    assign sel_R_DATA_TEMPR40  = (RAM_DEPTH > 32'h5000) ? int_R_DATA_TEMPR40  : 32'b0;
    assign sel_R_DATA_TEMPR41  = (RAM_DEPTH > 32'h5200) ? int_R_DATA_TEMPR41  : 32'b0;
    assign sel_R_DATA_TEMPR42  = (RAM_DEPTH > 32'h5400) ? int_R_DATA_TEMPR42  : 32'b0;
    assign sel_R_DATA_TEMPR43  = (RAM_DEPTH > 32'h5600) ? int_R_DATA_TEMPR43  : 32'b0;
    assign sel_R_DATA_TEMPR44  = (RAM_DEPTH > 32'h5800) ? int_R_DATA_TEMPR44  : 32'b0;
    assign sel_R_DATA_TEMPR45  = (RAM_DEPTH > 32'h5A00) ? int_R_DATA_TEMPR45  : 32'b0;
    assign sel_R_DATA_TEMPR46  = (RAM_DEPTH > 32'h5C00) ? int_R_DATA_TEMPR46  : 32'b0;
    assign sel_R_DATA_TEMPR47  = (RAM_DEPTH > 32'h5E00) ? int_R_DATA_TEMPR47  : 32'b0;
    assign sel_R_DATA_TEMPR48  = (RAM_DEPTH > 32'h6000) ? int_R_DATA_TEMPR48  : 32'b0;
    assign sel_R_DATA_TEMPR49  = (RAM_DEPTH > 32'h6200) ? int_R_DATA_TEMPR49  : 32'b0;
    assign sel_R_DATA_TEMPR50  = (RAM_DEPTH > 32'h6400) ? int_R_DATA_TEMPR50  : 32'b0;
    assign sel_R_DATA_TEMPR51  = (RAM_DEPTH > 32'h6600) ? int_R_DATA_TEMPR51  : 32'b0;
    assign sel_R_DATA_TEMPR52  = (RAM_DEPTH > 32'h6800) ? int_R_DATA_TEMPR52  : 32'b0;
    assign sel_R_DATA_TEMPR53  = (RAM_DEPTH > 32'h6A00) ? int_R_DATA_TEMPR53  : 32'b0;
    assign sel_R_DATA_TEMPR54  = (RAM_DEPTH > 32'h6C00) ? int_R_DATA_TEMPR54  : 32'b0;
    assign sel_R_DATA_TEMPR55  = (RAM_DEPTH > 32'h6E00) ? int_R_DATA_TEMPR55  : 32'b0;
    assign sel_R_DATA_TEMPR56  = (RAM_DEPTH > 32'h7000) ? int_R_DATA_TEMPR56  : 32'b0;
    assign sel_R_DATA_TEMPR57  = (RAM_DEPTH > 32'h7200) ? int_R_DATA_TEMPR57  : 32'b0;
    assign sel_R_DATA_TEMPR58  = (RAM_DEPTH > 32'h7400) ? int_R_DATA_TEMPR58  : 32'b0;
    assign sel_R_DATA_TEMPR59  = (RAM_DEPTH > 32'h7600) ? int_R_DATA_TEMPR59  : 32'b0;
    assign sel_R_DATA_TEMPR60  = (RAM_DEPTH > 32'h7800) ? int_R_DATA_TEMPR60  : 32'b0;
    assign sel_R_DATA_TEMPR61  = (RAM_DEPTH > 32'h7A00) ? int_R_DATA_TEMPR61  : 32'b0;
    assign sel_R_DATA_TEMPR62  = (RAM_DEPTH > 32'h7C00) ? int_R_DATA_TEMPR62  : 32'b0;
    assign sel_R_DATA_TEMPR63  = (RAM_DEPTH > 32'h7E00) ? int_R_DATA_TEMPR63  : 32'b0;
    assign sel_R_DATA_TEMPR64  = (RAM_DEPTH > 32'h8000) ? int_R_DATA_TEMPR64  : 32'b0;
    assign sel_R_DATA_TEMPR65  = (RAM_DEPTH > 32'h8200) ? int_R_DATA_TEMPR65  : 32'b0;
    assign sel_R_DATA_TEMPR66  = (RAM_DEPTH > 32'h8400) ? int_R_DATA_TEMPR66  : 32'b0;
    assign sel_R_DATA_TEMPR67  = (RAM_DEPTH > 32'h8600) ? int_R_DATA_TEMPR67  : 32'b0;
    assign sel_R_DATA_TEMPR68  = (RAM_DEPTH > 32'h8800) ? int_R_DATA_TEMPR68  : 32'b0;
    assign sel_R_DATA_TEMPR69  = (RAM_DEPTH > 32'h8A00) ? int_R_DATA_TEMPR69  : 32'b0;
    assign sel_R_DATA_TEMPR70  = (RAM_DEPTH > 32'h8C00) ? int_R_DATA_TEMPR70  : 32'b0;
    assign sel_R_DATA_TEMPR71  = (RAM_DEPTH > 32'h8E00) ? int_R_DATA_TEMPR71  : 32'b0;
    assign sel_R_DATA_TEMPR72  = (RAM_DEPTH > 32'h9000) ? int_R_DATA_TEMPR72  : 32'b0;
    assign sel_R_DATA_TEMPR73  = (RAM_DEPTH > 32'h9200) ? int_R_DATA_TEMPR73  : 32'b0;
    assign sel_R_DATA_TEMPR74  = (RAM_DEPTH > 32'h9400) ? int_R_DATA_TEMPR74  : 32'b0;
    assign sel_R_DATA_TEMPR75  = (RAM_DEPTH > 32'h9600) ? int_R_DATA_TEMPR75  : 32'b0;
    assign sel_R_DATA_TEMPR76  = (RAM_DEPTH > 32'h9800) ? int_R_DATA_TEMPR76  : 32'b0;
    assign sel_R_DATA_TEMPR77  = (RAM_DEPTH > 32'h9A00) ? int_R_DATA_TEMPR77  : 32'b0;
    assign sel_R_DATA_TEMPR78  = (RAM_DEPTH > 32'h9C00) ? int_R_DATA_TEMPR78  : 32'b0;
    assign sel_R_DATA_TEMPR79  = (RAM_DEPTH > 32'h9E00) ? int_R_DATA_TEMPR79  : 32'b0;
    assign sel_R_DATA_TEMPR80  = (RAM_DEPTH > 32'hA000) ? int_R_DATA_TEMPR80  : 32'b0;
    assign sel_R_DATA_TEMPR81  = (RAM_DEPTH > 32'hA200) ? int_R_DATA_TEMPR81  : 32'b0;
    assign sel_R_DATA_TEMPR82  = (RAM_DEPTH > 32'hA400) ? int_R_DATA_TEMPR82  : 32'b0;
    assign sel_R_DATA_TEMPR83  = (RAM_DEPTH > 32'hA600) ? int_R_DATA_TEMPR83  : 32'b0;
    assign sel_R_DATA_TEMPR84  = (RAM_DEPTH > 32'hA800) ? int_R_DATA_TEMPR84  : 32'b0;
    assign sel_R_DATA_TEMPR85  = (RAM_DEPTH > 32'hAA00) ? int_R_DATA_TEMPR85  : 32'b0;
    assign sel_R_DATA_TEMPR86  = (RAM_DEPTH > 32'hAC00) ? int_R_DATA_TEMPR86  : 32'b0;
    assign sel_R_DATA_TEMPR87  = (RAM_DEPTH > 32'hAE00) ? int_R_DATA_TEMPR87  : 32'b0;
    assign sel_R_DATA_TEMPR88  = (RAM_DEPTH > 32'hB000) ? int_R_DATA_TEMPR88  : 32'b0;
    assign sel_R_DATA_TEMPR89  = (RAM_DEPTH > 32'hB200) ? int_R_DATA_TEMPR89  : 32'b0;
    assign sel_R_DATA_TEMPR90  = (RAM_DEPTH > 32'hB400) ? int_R_DATA_TEMPR90  : 32'b0;
    assign sel_R_DATA_TEMPR91  = (RAM_DEPTH > 32'hB600) ? int_R_DATA_TEMPR91  : 32'b0;
    assign sel_R_DATA_TEMPR92  = (RAM_DEPTH > 32'hB800) ? int_R_DATA_TEMPR92  : 32'b0;
    assign sel_R_DATA_TEMPR93  = (RAM_DEPTH > 32'hBA00) ? int_R_DATA_TEMPR93  : 32'b0;
    assign sel_R_DATA_TEMPR94  = (RAM_DEPTH > 32'hBC00) ? int_R_DATA_TEMPR94  : 32'b0;
    assign sel_R_DATA_TEMPR95  = (RAM_DEPTH > 32'hBE00) ? int_R_DATA_TEMPR95  : 32'b0;
    assign sel_R_DATA_TEMPR96  = (RAM_DEPTH > 32'hC000) ? int_R_DATA_TEMPR96  : 32'b0;
    assign sel_R_DATA_TEMPR97  = (RAM_DEPTH > 32'hC200) ? int_R_DATA_TEMPR97  : 32'b0;
    assign sel_R_DATA_TEMPR98  = (RAM_DEPTH > 32'hC400) ? int_R_DATA_TEMPR98  : 32'b0;
    assign sel_R_DATA_TEMPR99  = (RAM_DEPTH > 32'hC600) ? int_R_DATA_TEMPR99  : 32'b0;
    assign sel_R_DATA_TEMPR100 = (RAM_DEPTH > 32'hC800) ? int_R_DATA_TEMPR100 : 32'b0;
    assign sel_R_DATA_TEMPR101 = (RAM_DEPTH > 32'hCA00) ? int_R_DATA_TEMPR101 : 32'b0;
    assign sel_R_DATA_TEMPR102 = (RAM_DEPTH > 32'hCC00) ? int_R_DATA_TEMPR102 : 32'b0;
    assign sel_R_DATA_TEMPR103 = (RAM_DEPTH > 32'hCE00) ? int_R_DATA_TEMPR103 : 32'b0;
    assign sel_R_DATA_TEMPR104 = (RAM_DEPTH > 32'hD000) ? int_R_DATA_TEMPR104 : 32'b0;
    assign sel_R_DATA_TEMPR105 = (RAM_DEPTH > 32'hD200) ? int_R_DATA_TEMPR105 : 32'b0;
    assign sel_R_DATA_TEMPR106 = (RAM_DEPTH > 32'hD400) ? int_R_DATA_TEMPR106 : 32'b0;
    assign sel_R_DATA_TEMPR107 = (RAM_DEPTH > 32'hD600) ? int_R_DATA_TEMPR107 : 32'b0;
    assign sel_R_DATA_TEMPR108 = (RAM_DEPTH > 32'hD800) ? int_R_DATA_TEMPR108 : 32'b0;
    assign sel_R_DATA_TEMPR109 = (RAM_DEPTH > 32'hDA00) ? int_R_DATA_TEMPR109 : 32'b0;
    assign sel_R_DATA_TEMPR110 = (RAM_DEPTH > 32'hDC00) ? int_R_DATA_TEMPR110 : 32'b0;
    assign sel_R_DATA_TEMPR111 = (RAM_DEPTH > 32'hDE00) ? int_R_DATA_TEMPR111 : 32'b0;
    assign sel_R_DATA_TEMPR112 = (RAM_DEPTH > 32'hE000) ? int_R_DATA_TEMPR112 : 32'b0;
    assign sel_R_DATA_TEMPR113 = (RAM_DEPTH > 32'hE200) ? int_R_DATA_TEMPR113 : 32'b0;
    assign sel_R_DATA_TEMPR114 = (RAM_DEPTH > 32'hE400) ? int_R_DATA_TEMPR114 : 32'b0;
    assign sel_R_DATA_TEMPR115 = (RAM_DEPTH > 32'hE600) ? int_R_DATA_TEMPR115 : 32'b0;
    assign sel_R_DATA_TEMPR116 = (RAM_DEPTH > 32'hE800) ? int_R_DATA_TEMPR116 : 32'b0;
    assign sel_R_DATA_TEMPR117 = (RAM_DEPTH > 32'hEA00) ? int_R_DATA_TEMPR117 : 32'b0;
    assign sel_R_DATA_TEMPR118 = (RAM_DEPTH > 32'hEC00) ? int_R_DATA_TEMPR118 : 32'b0;
    assign sel_R_DATA_TEMPR119 = (RAM_DEPTH > 32'hEE00) ? int_R_DATA_TEMPR119 : 32'b0;
    assign sel_R_DATA_TEMPR120 = (RAM_DEPTH > 32'hF000) ? int_R_DATA_TEMPR120 : 32'b0;
    assign sel_R_DATA_TEMPR121 = (RAM_DEPTH > 32'hF200) ? int_R_DATA_TEMPR121 : 32'b0;
    assign sel_R_DATA_TEMPR122 = (RAM_DEPTH > 32'hF400) ? int_R_DATA_TEMPR122 : 32'b0;
    assign sel_R_DATA_TEMPR123 = (RAM_DEPTH > 32'hF600) ? int_R_DATA_TEMPR123 : 32'b0;
    assign sel_R_DATA_TEMPR124 = (RAM_DEPTH > 32'hF800) ? int_R_DATA_TEMPR124 : 32'b0;
    assign sel_R_DATA_TEMPR125 = (RAM_DEPTH > 32'hFA00) ? int_R_DATA_TEMPR125 : 32'b0;
    assign sel_R_DATA_TEMPR126 = (RAM_DEPTH > 32'hFC00) ? int_R_DATA_TEMPR126 : 32'b0;
    assign sel_R_DATA_TEMPR127 = (RAM_DEPTH > 32'hFE00) ? int_R_DATA_TEMPR127 : 32'b0;
	
    assign sel_SB_CORRECT_NG[0  ] = (RAM_DEPTH > 32'h0   ) ? int_SB_CORRECT_NG[0  ] : 1'b0;
    assign sel_SB_CORRECT_NG[1  ] = (RAM_DEPTH > 32'h200 ) ? int_SB_CORRECT_NG[1  ] : 1'b0;
    assign sel_SB_CORRECT_NG[2  ] = (RAM_DEPTH > 32'h400 ) ? int_SB_CORRECT_NG[2  ] : 1'b0;
    assign sel_SB_CORRECT_NG[3  ] = (RAM_DEPTH > 32'h600 ) ? int_SB_CORRECT_NG[3  ] : 1'b0;
    assign sel_SB_CORRECT_NG[4  ] = (RAM_DEPTH > 32'h800 ) ? int_SB_CORRECT_NG[4  ] : 1'b0;
    assign sel_SB_CORRECT_NG[5  ] = (RAM_DEPTH > 32'hA00 ) ? int_SB_CORRECT_NG[5  ] : 1'b0;
    assign sel_SB_CORRECT_NG[6  ] = (RAM_DEPTH > 32'hC00 ) ? int_SB_CORRECT_NG[6  ] : 1'b0;
    assign sel_SB_CORRECT_NG[7  ] = (RAM_DEPTH > 32'hE00 ) ? int_SB_CORRECT_NG[7  ] : 1'b0;
    assign sel_SB_CORRECT_NG[8  ] = (RAM_DEPTH > 32'h1000) ? int_SB_CORRECT_NG[8  ] : 1'b0;
    assign sel_SB_CORRECT_NG[9  ] = (RAM_DEPTH > 32'h1200) ? int_SB_CORRECT_NG[9  ] : 1'b0;
    assign sel_SB_CORRECT_NG[10 ] = (RAM_DEPTH > 32'h1400) ? int_SB_CORRECT_NG[10 ] : 1'b0;
    assign sel_SB_CORRECT_NG[11 ] = (RAM_DEPTH > 32'h1600) ? int_SB_CORRECT_NG[11 ] : 1'b0;
    assign sel_SB_CORRECT_NG[12 ] = (RAM_DEPTH > 32'h1800) ? int_SB_CORRECT_NG[12 ] : 1'b0;
    assign sel_SB_CORRECT_NG[13 ] = (RAM_DEPTH > 32'h1A00) ? int_SB_CORRECT_NG[13 ] : 1'b0;
    assign sel_SB_CORRECT_NG[14 ] = (RAM_DEPTH > 32'h1C00) ? int_SB_CORRECT_NG[14 ] : 1'b0;
    assign sel_SB_CORRECT_NG[15 ] = (RAM_DEPTH > 32'h1E00) ? int_SB_CORRECT_NG[15 ] : 1'b0;
    assign sel_SB_CORRECT_NG[16 ] = (RAM_DEPTH > 32'h2000) ? int_SB_CORRECT_NG[16 ] : 1'b0;
    assign sel_SB_CORRECT_NG[17 ] = (RAM_DEPTH > 32'h2200) ? int_SB_CORRECT_NG[17 ] : 1'b0;
    assign sel_SB_CORRECT_NG[18 ] = (RAM_DEPTH > 32'h2400) ? int_SB_CORRECT_NG[18 ] : 1'b0;
    assign sel_SB_CORRECT_NG[19 ] = (RAM_DEPTH > 32'h2600) ? int_SB_CORRECT_NG[19 ] : 1'b0;
    assign sel_SB_CORRECT_NG[20 ] = (RAM_DEPTH > 32'h2800) ? int_SB_CORRECT_NG[20 ] : 1'b0;
    assign sel_SB_CORRECT_NG[21 ] = (RAM_DEPTH > 32'h2A00) ? int_SB_CORRECT_NG[21 ] : 1'b0;
    assign sel_SB_CORRECT_NG[22 ] = (RAM_DEPTH > 32'h2C00) ? int_SB_CORRECT_NG[22 ] : 1'b0;
    assign sel_SB_CORRECT_NG[23 ] = (RAM_DEPTH > 32'h2E00) ? int_SB_CORRECT_NG[23 ] : 1'b0;
    assign sel_SB_CORRECT_NG[24 ] = (RAM_DEPTH > 32'h3000) ? int_SB_CORRECT_NG[24 ] : 1'b0;
    assign sel_SB_CORRECT_NG[25 ] = (RAM_DEPTH > 32'h3200) ? int_SB_CORRECT_NG[25 ] : 1'b0;
    assign sel_SB_CORRECT_NG[26 ] = (RAM_DEPTH > 32'h3400) ? int_SB_CORRECT_NG[26 ] : 1'b0;
    assign sel_SB_CORRECT_NG[27 ] = (RAM_DEPTH > 32'h3600) ? int_SB_CORRECT_NG[27 ] : 1'b0;
    assign sel_SB_CORRECT_NG[28 ] = (RAM_DEPTH > 32'h3800) ? int_SB_CORRECT_NG[28 ] : 1'b0;
    assign sel_SB_CORRECT_NG[29 ] = (RAM_DEPTH > 32'h3A00) ? int_SB_CORRECT_NG[29 ] : 1'b0;
    assign sel_SB_CORRECT_NG[30 ] = (RAM_DEPTH > 32'h3C00) ? int_SB_CORRECT_NG[30 ] : 1'b0;
    assign sel_SB_CORRECT_NG[31 ] = (RAM_DEPTH > 32'h3E00) ? int_SB_CORRECT_NG[31 ] : 1'b0;
    assign sel_SB_CORRECT_NG[32 ] = (RAM_DEPTH > 32'h4000) ? int_SB_CORRECT_NG[32 ] : 1'b0;
    assign sel_SB_CORRECT_NG[33 ] = (RAM_DEPTH > 32'h4200) ? int_SB_CORRECT_NG[33 ] : 1'b0;
    assign sel_SB_CORRECT_NG[34 ] = (RAM_DEPTH > 32'h4400) ? int_SB_CORRECT_NG[34 ] : 1'b0;
    assign sel_SB_CORRECT_NG[35 ] = (RAM_DEPTH > 32'h4600) ? int_SB_CORRECT_NG[35 ] : 1'b0;
    assign sel_SB_CORRECT_NG[36 ] = (RAM_DEPTH > 32'h4800) ? int_SB_CORRECT_NG[36 ] : 1'b0;
    assign sel_SB_CORRECT_NG[37 ] = (RAM_DEPTH > 32'h4A00) ? int_SB_CORRECT_NG[37 ] : 1'b0;
    assign sel_SB_CORRECT_NG[38 ] = (RAM_DEPTH > 32'h4C00) ? int_SB_CORRECT_NG[38 ] : 1'b0;
    assign sel_SB_CORRECT_NG[39 ] = (RAM_DEPTH > 32'h4E00) ? int_SB_CORRECT_NG[39 ] : 1'b0;
    assign sel_SB_CORRECT_NG[40 ] = (RAM_DEPTH > 32'h5000) ? int_SB_CORRECT_NG[40 ] : 1'b0;
    assign sel_SB_CORRECT_NG[41 ] = (RAM_DEPTH > 32'h5200) ? int_SB_CORRECT_NG[41 ] : 1'b0;
    assign sel_SB_CORRECT_NG[42 ] = (RAM_DEPTH > 32'h5400) ? int_SB_CORRECT_NG[42 ] : 1'b0;
    assign sel_SB_CORRECT_NG[43 ] = (RAM_DEPTH > 32'h5600) ? int_SB_CORRECT_NG[43 ] : 1'b0;
    assign sel_SB_CORRECT_NG[44 ] = (RAM_DEPTH > 32'h5800) ? int_SB_CORRECT_NG[44 ] : 1'b0;
    assign sel_SB_CORRECT_NG[45 ] = (RAM_DEPTH > 32'h5A00) ? int_SB_CORRECT_NG[45 ] : 1'b0;
    assign sel_SB_CORRECT_NG[46 ] = (RAM_DEPTH > 32'h5C00) ? int_SB_CORRECT_NG[46 ] : 1'b0;
    assign sel_SB_CORRECT_NG[47 ] = (RAM_DEPTH > 32'h5E00) ? int_SB_CORRECT_NG[47 ] : 1'b0;
    assign sel_SB_CORRECT_NG[48 ] = (RAM_DEPTH > 32'h6000) ? int_SB_CORRECT_NG[48 ] : 1'b0;
    assign sel_SB_CORRECT_NG[49 ] = (RAM_DEPTH > 32'h6200) ? int_SB_CORRECT_NG[49 ] : 1'b0;
    assign sel_SB_CORRECT_NG[50 ] = (RAM_DEPTH > 32'h6400) ? int_SB_CORRECT_NG[50 ] : 1'b0;
    assign sel_SB_CORRECT_NG[51 ] = (RAM_DEPTH > 32'h6600) ? int_SB_CORRECT_NG[51 ] : 1'b0;
    assign sel_SB_CORRECT_NG[52 ] = (RAM_DEPTH > 32'h6800) ? int_SB_CORRECT_NG[52 ] : 1'b0;
    assign sel_SB_CORRECT_NG[53 ] = (RAM_DEPTH > 32'h6A00) ? int_SB_CORRECT_NG[53 ] : 1'b0;
    assign sel_SB_CORRECT_NG[54 ] = (RAM_DEPTH > 32'h6C00) ? int_SB_CORRECT_NG[54 ] : 1'b0;
    assign sel_SB_CORRECT_NG[55 ] = (RAM_DEPTH > 32'h6E00) ? int_SB_CORRECT_NG[55 ] : 1'b0;
    assign sel_SB_CORRECT_NG[56 ] = (RAM_DEPTH > 32'h7000) ? int_SB_CORRECT_NG[56 ] : 1'b0;
    assign sel_SB_CORRECT_NG[57 ] = (RAM_DEPTH > 32'h7200) ? int_SB_CORRECT_NG[57 ] : 1'b0;
    assign sel_SB_CORRECT_NG[58 ] = (RAM_DEPTH > 32'h7400) ? int_SB_CORRECT_NG[58 ] : 1'b0;
    assign sel_SB_CORRECT_NG[59 ] = (RAM_DEPTH > 32'h7600) ? int_SB_CORRECT_NG[59 ] : 1'b0;
    assign sel_SB_CORRECT_NG[60 ] = (RAM_DEPTH > 32'h7800) ? int_SB_CORRECT_NG[60 ] : 1'b0;
    assign sel_SB_CORRECT_NG[61 ] = (RAM_DEPTH > 32'h7A00) ? int_SB_CORRECT_NG[61 ] : 1'b0;
    assign sel_SB_CORRECT_NG[62 ] = (RAM_DEPTH > 32'h7C00) ? int_SB_CORRECT_NG[62 ] : 1'b0;
    assign sel_SB_CORRECT_NG[63 ] = (RAM_DEPTH > 32'h7E00) ? int_SB_CORRECT_NG[63 ] : 1'b0;
    assign sel_SB_CORRECT_NG[64 ] = (RAM_DEPTH > 32'h8000) ? int_SB_CORRECT_NG[64 ] : 1'b0;
    assign sel_SB_CORRECT_NG[65 ] = (RAM_DEPTH > 32'h8200) ? int_SB_CORRECT_NG[65 ] : 1'b0;
    assign sel_SB_CORRECT_NG[66 ] = (RAM_DEPTH > 32'h8400) ? int_SB_CORRECT_NG[66 ] : 1'b0;
    assign sel_SB_CORRECT_NG[67 ] = (RAM_DEPTH > 32'h8600) ? int_SB_CORRECT_NG[67 ] : 1'b0;
    assign sel_SB_CORRECT_NG[68 ] = (RAM_DEPTH > 32'h8800) ? int_SB_CORRECT_NG[68 ] : 1'b0;
    assign sel_SB_CORRECT_NG[69 ] = (RAM_DEPTH > 32'h8A00) ? int_SB_CORRECT_NG[69 ] : 1'b0;
    assign sel_SB_CORRECT_NG[70 ] = (RAM_DEPTH > 32'h8C00) ? int_SB_CORRECT_NG[70 ] : 1'b0;
    assign sel_SB_CORRECT_NG[71 ] = (RAM_DEPTH > 32'h8E00) ? int_SB_CORRECT_NG[71 ] : 1'b0;
    assign sel_SB_CORRECT_NG[72 ] = (RAM_DEPTH > 32'h9000) ? int_SB_CORRECT_NG[72 ] : 1'b0;
    assign sel_SB_CORRECT_NG[73 ] = (RAM_DEPTH > 32'h9200) ? int_SB_CORRECT_NG[73 ] : 1'b0;
    assign sel_SB_CORRECT_NG[74 ] = (RAM_DEPTH > 32'h9400) ? int_SB_CORRECT_NG[74 ] : 1'b0;
    assign sel_SB_CORRECT_NG[75 ] = (RAM_DEPTH > 32'h9600) ? int_SB_CORRECT_NG[75 ] : 1'b0;
    assign sel_SB_CORRECT_NG[76 ] = (RAM_DEPTH > 32'h9800) ? int_SB_CORRECT_NG[76 ] : 1'b0;
    assign sel_SB_CORRECT_NG[77 ] = (RAM_DEPTH > 32'h9A00) ? int_SB_CORRECT_NG[77 ] : 1'b0;
    assign sel_SB_CORRECT_NG[78 ] = (RAM_DEPTH > 32'h9C00) ? int_SB_CORRECT_NG[78 ] : 1'b0;
    assign sel_SB_CORRECT_NG[79 ] = (RAM_DEPTH > 32'h9E00) ? int_SB_CORRECT_NG[79 ] : 1'b0;
    assign sel_SB_CORRECT_NG[80 ] = (RAM_DEPTH > 32'hA000) ? int_SB_CORRECT_NG[80 ] : 1'b0;
    assign sel_SB_CORRECT_NG[81 ] = (RAM_DEPTH > 32'hA200) ? int_SB_CORRECT_NG[81 ] : 1'b0;
    assign sel_SB_CORRECT_NG[82 ] = (RAM_DEPTH > 32'hA400) ? int_SB_CORRECT_NG[82 ] : 1'b0;
    assign sel_SB_CORRECT_NG[83 ] = (RAM_DEPTH > 32'hA600) ? int_SB_CORRECT_NG[83 ] : 1'b0;
    assign sel_SB_CORRECT_NG[84 ] = (RAM_DEPTH > 32'hA800) ? int_SB_CORRECT_NG[84 ] : 1'b0;
    assign sel_SB_CORRECT_NG[85 ] = (RAM_DEPTH > 32'hAA00) ? int_SB_CORRECT_NG[85 ] : 1'b0;
    assign sel_SB_CORRECT_NG[86 ] = (RAM_DEPTH > 32'hAC00) ? int_SB_CORRECT_NG[86 ] : 1'b0;
    assign sel_SB_CORRECT_NG[87 ] = (RAM_DEPTH > 32'hAE00) ? int_SB_CORRECT_NG[87 ] : 1'b0;
    assign sel_SB_CORRECT_NG[88 ] = (RAM_DEPTH > 32'hB000) ? int_SB_CORRECT_NG[88 ] : 1'b0;
    assign sel_SB_CORRECT_NG[89 ] = (RAM_DEPTH > 32'hB200) ? int_SB_CORRECT_NG[89 ] : 1'b0;
    assign sel_SB_CORRECT_NG[90 ] = (RAM_DEPTH > 32'hB400) ? int_SB_CORRECT_NG[90 ] : 1'b0;
    assign sel_SB_CORRECT_NG[91 ] = (RAM_DEPTH > 32'hB600) ? int_SB_CORRECT_NG[91 ] : 1'b0;
    assign sel_SB_CORRECT_NG[92 ] = (RAM_DEPTH > 32'hB800) ? int_SB_CORRECT_NG[92 ] : 1'b0;
    assign sel_SB_CORRECT_NG[93 ] = (RAM_DEPTH > 32'hBA00) ? int_SB_CORRECT_NG[93 ] : 1'b0;
    assign sel_SB_CORRECT_NG[94 ] = (RAM_DEPTH > 32'hBC00) ? int_SB_CORRECT_NG[94 ] : 1'b0;
    assign sel_SB_CORRECT_NG[95 ] = (RAM_DEPTH > 32'hBE00) ? int_SB_CORRECT_NG[95 ] : 1'b0;
    assign sel_SB_CORRECT_NG[96 ] = (RAM_DEPTH > 32'hC000) ? int_SB_CORRECT_NG[96 ] : 1'b0;
    assign sel_SB_CORRECT_NG[97 ] = (RAM_DEPTH > 32'hC200) ? int_SB_CORRECT_NG[97 ] : 1'b0;
    assign sel_SB_CORRECT_NG[98 ] = (RAM_DEPTH > 32'hC400) ? int_SB_CORRECT_NG[98 ] : 1'b0;
    assign sel_SB_CORRECT_NG[99 ] = (RAM_DEPTH > 32'hC600) ? int_SB_CORRECT_NG[99 ] : 1'b0;
    assign sel_SB_CORRECT_NG[100] = (RAM_DEPTH > 32'hC800) ? int_SB_CORRECT_NG[100] : 1'b0;
    assign sel_SB_CORRECT_NG[101] = (RAM_DEPTH > 32'hCA00) ? int_SB_CORRECT_NG[101] : 1'b0;
    assign sel_SB_CORRECT_NG[102] = (RAM_DEPTH > 32'hCC00) ? int_SB_CORRECT_NG[102] : 1'b0;
    assign sel_SB_CORRECT_NG[103] = (RAM_DEPTH > 32'hCE00) ? int_SB_CORRECT_NG[103] : 1'b0;
    assign sel_SB_CORRECT_NG[104] = (RAM_DEPTH > 32'hD000) ? int_SB_CORRECT_NG[104] : 1'b0;
    assign sel_SB_CORRECT_NG[105] = (RAM_DEPTH > 32'hD200) ? int_SB_CORRECT_NG[105] : 1'b0;
    assign sel_SB_CORRECT_NG[106] = (RAM_DEPTH > 32'hD400) ? int_SB_CORRECT_NG[106] : 1'b0;
    assign sel_SB_CORRECT_NG[107] = (RAM_DEPTH > 32'hD600) ? int_SB_CORRECT_NG[107] : 1'b0;
    assign sel_SB_CORRECT_NG[108] = (RAM_DEPTH > 32'hD800) ? int_SB_CORRECT_NG[108] : 1'b0;
    assign sel_SB_CORRECT_NG[109] = (RAM_DEPTH > 32'hDA00) ? int_SB_CORRECT_NG[109] : 1'b0;
    assign sel_SB_CORRECT_NG[110] = (RAM_DEPTH > 32'hDC00) ? int_SB_CORRECT_NG[110] : 1'b0;
    assign sel_SB_CORRECT_NG[111] = (RAM_DEPTH > 32'hDE00) ? int_SB_CORRECT_NG[111] : 1'b0;
    assign sel_SB_CORRECT_NG[112] = (RAM_DEPTH > 32'hE000) ? int_SB_CORRECT_NG[112] : 1'b0;
    assign sel_SB_CORRECT_NG[113] = (RAM_DEPTH > 32'hE200) ? int_SB_CORRECT_NG[113] : 1'b0;
    assign sel_SB_CORRECT_NG[114] = (RAM_DEPTH > 32'hE400) ? int_SB_CORRECT_NG[114] : 1'b0;
    assign sel_SB_CORRECT_NG[115] = (RAM_DEPTH > 32'hE600) ? int_SB_CORRECT_NG[115] : 1'b0;
    assign sel_SB_CORRECT_NG[116] = (RAM_DEPTH > 32'hE800) ? int_SB_CORRECT_NG[116] : 1'b0;
    assign sel_SB_CORRECT_NG[117] = (RAM_DEPTH > 32'hEA00) ? int_SB_CORRECT_NG[117] : 1'b0;
    assign sel_SB_CORRECT_NG[118] = (RAM_DEPTH > 32'hEC00) ? int_SB_CORRECT_NG[118] : 1'b0;
    assign sel_SB_CORRECT_NG[119] = (RAM_DEPTH > 32'hEE00) ? int_SB_CORRECT_NG[119] : 1'b0;
    assign sel_SB_CORRECT_NG[120] = (RAM_DEPTH > 32'hF000) ? int_SB_CORRECT_NG[120] : 1'b0;
    assign sel_SB_CORRECT_NG[121] = (RAM_DEPTH > 32'hF200) ? int_SB_CORRECT_NG[121] : 1'b0;
    assign sel_SB_CORRECT_NG[122] = (RAM_DEPTH > 32'hF400) ? int_SB_CORRECT_NG[122] : 1'b0;
    assign sel_SB_CORRECT_NG[123] = (RAM_DEPTH > 32'hF600) ? int_SB_CORRECT_NG[123] : 1'b0;
    assign sel_SB_CORRECT_NG[124] = (RAM_DEPTH > 32'hF800) ? int_SB_CORRECT_NG[124] : 1'b0;
    assign sel_SB_CORRECT_NG[125] = (RAM_DEPTH > 32'hFA00) ? int_SB_CORRECT_NG[125] : 1'b0;
    assign sel_SB_CORRECT_NG[126] = (RAM_DEPTH > 32'hFC00) ? int_SB_CORRECT_NG[126] : 1'b0;
    assign sel_SB_CORRECT_NG[127] = (RAM_DEPTH > 32'hFE00) ? int_SB_CORRECT_NG[127] : 1'b0;
	
    assign sel_DB_DETECT_NG[0  ] = (RAM_DEPTH > 32'h0   ) ? int_DB_DETECT_NG[0  ] : 1'b0;
    assign sel_DB_DETECT_NG[1  ] = (RAM_DEPTH > 32'h200 ) ? int_DB_DETECT_NG[1  ] : 1'b0;
    assign sel_DB_DETECT_NG[2  ] = (RAM_DEPTH > 32'h400 ) ? int_DB_DETECT_NG[2  ] : 1'b0;
    assign sel_DB_DETECT_NG[3  ] = (RAM_DEPTH > 32'h600 ) ? int_DB_DETECT_NG[3  ] : 1'b0;
    assign sel_DB_DETECT_NG[4  ] = (RAM_DEPTH > 32'h800 ) ? int_DB_DETECT_NG[4  ] : 1'b0;
    assign sel_DB_DETECT_NG[5  ] = (RAM_DEPTH > 32'hA00 ) ? int_DB_DETECT_NG[5  ] : 1'b0;
    assign sel_DB_DETECT_NG[6  ] = (RAM_DEPTH > 32'hC00 ) ? int_DB_DETECT_NG[6  ] : 1'b0;
    assign sel_DB_DETECT_NG[7  ] = (RAM_DEPTH > 32'hE00 ) ? int_DB_DETECT_NG[7  ] : 1'b0;
    assign sel_DB_DETECT_NG[8  ] = (RAM_DEPTH > 32'h1000) ? int_DB_DETECT_NG[8  ] : 1'b0;
    assign sel_DB_DETECT_NG[9  ] = (RAM_DEPTH > 32'h1200) ? int_DB_DETECT_NG[9  ] : 1'b0;
    assign sel_DB_DETECT_NG[10 ] = (RAM_DEPTH > 32'h1400) ? int_DB_DETECT_NG[10 ] : 1'b0;
    assign sel_DB_DETECT_NG[11 ] = (RAM_DEPTH > 32'h1600) ? int_DB_DETECT_NG[11 ] : 1'b0;
    assign sel_DB_DETECT_NG[12 ] = (RAM_DEPTH > 32'h1800) ? int_DB_DETECT_NG[12 ] : 1'b0;
    assign sel_DB_DETECT_NG[13 ] = (RAM_DEPTH > 32'h1A00) ? int_DB_DETECT_NG[13 ] : 1'b0;
    assign sel_DB_DETECT_NG[14 ] = (RAM_DEPTH > 32'h1C00) ? int_DB_DETECT_NG[14 ] : 1'b0;
    assign sel_DB_DETECT_NG[15 ] = (RAM_DEPTH > 32'h1E00) ? int_DB_DETECT_NG[15 ] : 1'b0;
    assign sel_DB_DETECT_NG[16 ] = (RAM_DEPTH > 32'h2000) ? int_DB_DETECT_NG[16 ] : 1'b0;
    assign sel_DB_DETECT_NG[17 ] = (RAM_DEPTH > 32'h2200) ? int_DB_DETECT_NG[17 ] : 1'b0;
    assign sel_DB_DETECT_NG[18 ] = (RAM_DEPTH > 32'h2400) ? int_DB_DETECT_NG[18 ] : 1'b0;
    assign sel_DB_DETECT_NG[19 ] = (RAM_DEPTH > 32'h2600) ? int_DB_DETECT_NG[19 ] : 1'b0;
    assign sel_DB_DETECT_NG[20 ] = (RAM_DEPTH > 32'h2800) ? int_DB_DETECT_NG[20 ] : 1'b0;
    assign sel_DB_DETECT_NG[21 ] = (RAM_DEPTH > 32'h2A00) ? int_DB_DETECT_NG[21 ] : 1'b0;
    assign sel_DB_DETECT_NG[22 ] = (RAM_DEPTH > 32'h2C00) ? int_DB_DETECT_NG[22 ] : 1'b0;
    assign sel_DB_DETECT_NG[23 ] = (RAM_DEPTH > 32'h2E00) ? int_DB_DETECT_NG[23 ] : 1'b0;
    assign sel_DB_DETECT_NG[24 ] = (RAM_DEPTH > 32'h3000) ? int_DB_DETECT_NG[24 ] : 1'b0;
    assign sel_DB_DETECT_NG[25 ] = (RAM_DEPTH > 32'h3200) ? int_DB_DETECT_NG[25 ] : 1'b0;
    assign sel_DB_DETECT_NG[26 ] = (RAM_DEPTH > 32'h3400) ? int_DB_DETECT_NG[26 ] : 1'b0;
    assign sel_DB_DETECT_NG[27 ] = (RAM_DEPTH > 32'h3600) ? int_DB_DETECT_NG[27 ] : 1'b0;
    assign sel_DB_DETECT_NG[28 ] = (RAM_DEPTH > 32'h3800) ? int_DB_DETECT_NG[28 ] : 1'b0;
    assign sel_DB_DETECT_NG[29 ] = (RAM_DEPTH > 32'h3A00) ? int_DB_DETECT_NG[29 ] : 1'b0;
    assign sel_DB_DETECT_NG[30 ] = (RAM_DEPTH > 32'h3C00) ? int_DB_DETECT_NG[30 ] : 1'b0;
    assign sel_DB_DETECT_NG[31 ] = (RAM_DEPTH > 32'h3E00) ? int_DB_DETECT_NG[31 ] : 1'b0;
    assign sel_DB_DETECT_NG[32 ] = (RAM_DEPTH > 32'h4000) ? int_DB_DETECT_NG[32 ] : 1'b0;
    assign sel_DB_DETECT_NG[33 ] = (RAM_DEPTH > 32'h4200) ? int_DB_DETECT_NG[33 ] : 1'b0;
    assign sel_DB_DETECT_NG[34 ] = (RAM_DEPTH > 32'h4400) ? int_DB_DETECT_NG[34 ] : 1'b0;
    assign sel_DB_DETECT_NG[35 ] = (RAM_DEPTH > 32'h4600) ? int_DB_DETECT_NG[35 ] : 1'b0;
    assign sel_DB_DETECT_NG[36 ] = (RAM_DEPTH > 32'h4800) ? int_DB_DETECT_NG[36 ] : 1'b0;
    assign sel_DB_DETECT_NG[37 ] = (RAM_DEPTH > 32'h4A00) ? int_DB_DETECT_NG[37 ] : 1'b0;
    assign sel_DB_DETECT_NG[38 ] = (RAM_DEPTH > 32'h4C00) ? int_DB_DETECT_NG[38 ] : 1'b0;
    assign sel_DB_DETECT_NG[39 ] = (RAM_DEPTH > 32'h4E00) ? int_DB_DETECT_NG[39 ] : 1'b0;
    assign sel_DB_DETECT_NG[40 ] = (RAM_DEPTH > 32'h5000) ? int_DB_DETECT_NG[40 ] : 1'b0;
    assign sel_DB_DETECT_NG[41 ] = (RAM_DEPTH > 32'h5200) ? int_DB_DETECT_NG[41 ] : 1'b0;
    assign sel_DB_DETECT_NG[42 ] = (RAM_DEPTH > 32'h5400) ? int_DB_DETECT_NG[42 ] : 1'b0;
    assign sel_DB_DETECT_NG[43 ] = (RAM_DEPTH > 32'h5600) ? int_DB_DETECT_NG[43 ] : 1'b0;
    assign sel_DB_DETECT_NG[44 ] = (RAM_DEPTH > 32'h5800) ? int_DB_DETECT_NG[44 ] : 1'b0;
    assign sel_DB_DETECT_NG[45 ] = (RAM_DEPTH > 32'h5A00) ? int_DB_DETECT_NG[45 ] : 1'b0;
    assign sel_DB_DETECT_NG[46 ] = (RAM_DEPTH > 32'h5C00) ? int_DB_DETECT_NG[46 ] : 1'b0;
    assign sel_DB_DETECT_NG[47 ] = (RAM_DEPTH > 32'h5E00) ? int_DB_DETECT_NG[47 ] : 1'b0;
    assign sel_DB_DETECT_NG[48 ] = (RAM_DEPTH > 32'h6000) ? int_DB_DETECT_NG[48 ] : 1'b0;
    assign sel_DB_DETECT_NG[49 ] = (RAM_DEPTH > 32'h6200) ? int_DB_DETECT_NG[49 ] : 1'b0;
    assign sel_DB_DETECT_NG[50 ] = (RAM_DEPTH > 32'h6400) ? int_DB_DETECT_NG[50 ] : 1'b0;
    assign sel_DB_DETECT_NG[51 ] = (RAM_DEPTH > 32'h6600) ? int_DB_DETECT_NG[51 ] : 1'b0;
    assign sel_DB_DETECT_NG[52 ] = (RAM_DEPTH > 32'h6800) ? int_DB_DETECT_NG[52 ] : 1'b0;
    assign sel_DB_DETECT_NG[53 ] = (RAM_DEPTH > 32'h6A00) ? int_DB_DETECT_NG[53 ] : 1'b0;
    assign sel_DB_DETECT_NG[54 ] = (RAM_DEPTH > 32'h6C00) ? int_DB_DETECT_NG[54 ] : 1'b0;
    assign sel_DB_DETECT_NG[55 ] = (RAM_DEPTH > 32'h6E00) ? int_DB_DETECT_NG[55 ] : 1'b0;
    assign sel_DB_DETECT_NG[56 ] = (RAM_DEPTH > 32'h7000) ? int_DB_DETECT_NG[56 ] : 1'b0;
    assign sel_DB_DETECT_NG[57 ] = (RAM_DEPTH > 32'h7200) ? int_DB_DETECT_NG[57 ] : 1'b0;
    assign sel_DB_DETECT_NG[58 ] = (RAM_DEPTH > 32'h7400) ? int_DB_DETECT_NG[58 ] : 1'b0;
    assign sel_DB_DETECT_NG[59 ] = (RAM_DEPTH > 32'h7600) ? int_DB_DETECT_NG[59 ] : 1'b0;
    assign sel_DB_DETECT_NG[60 ] = (RAM_DEPTH > 32'h7800) ? int_DB_DETECT_NG[60 ] : 1'b0;
    assign sel_DB_DETECT_NG[61 ] = (RAM_DEPTH > 32'h7A00) ? int_DB_DETECT_NG[61 ] : 1'b0;
    assign sel_DB_DETECT_NG[62 ] = (RAM_DEPTH > 32'h7C00) ? int_DB_DETECT_NG[62 ] : 1'b0;
    assign sel_DB_DETECT_NG[63 ] = (RAM_DEPTH > 32'h7E00) ? int_DB_DETECT_NG[63 ] : 1'b0;
    assign sel_DB_DETECT_NG[64 ] = (RAM_DEPTH > 32'h8000) ? int_DB_DETECT_NG[64 ] : 1'b0;
    assign sel_DB_DETECT_NG[65 ] = (RAM_DEPTH > 32'h8200) ? int_DB_DETECT_NG[65 ] : 1'b0;
    assign sel_DB_DETECT_NG[66 ] = (RAM_DEPTH > 32'h8400) ? int_DB_DETECT_NG[66 ] : 1'b0;
    assign sel_DB_DETECT_NG[67 ] = (RAM_DEPTH > 32'h8600) ? int_DB_DETECT_NG[67 ] : 1'b0;
    assign sel_DB_DETECT_NG[68 ] = (RAM_DEPTH > 32'h8800) ? int_DB_DETECT_NG[68 ] : 1'b0;
    assign sel_DB_DETECT_NG[69 ] = (RAM_DEPTH > 32'h8A00) ? int_DB_DETECT_NG[69 ] : 1'b0;
    assign sel_DB_DETECT_NG[70 ] = (RAM_DEPTH > 32'h8C00) ? int_DB_DETECT_NG[70 ] : 1'b0;
    assign sel_DB_DETECT_NG[71 ] = (RAM_DEPTH > 32'h8E00) ? int_DB_DETECT_NG[71 ] : 1'b0;
    assign sel_DB_DETECT_NG[72 ] = (RAM_DEPTH > 32'h9000) ? int_DB_DETECT_NG[72 ] : 1'b0;
    assign sel_DB_DETECT_NG[73 ] = (RAM_DEPTH > 32'h9200) ? int_DB_DETECT_NG[73 ] : 1'b0;
    assign sel_DB_DETECT_NG[74 ] = (RAM_DEPTH > 32'h9400) ? int_DB_DETECT_NG[74 ] : 1'b0;
    assign sel_DB_DETECT_NG[75 ] = (RAM_DEPTH > 32'h9600) ? int_DB_DETECT_NG[75 ] : 1'b0;
    assign sel_DB_DETECT_NG[76 ] = (RAM_DEPTH > 32'h9800) ? int_DB_DETECT_NG[76 ] : 1'b0;
    assign sel_DB_DETECT_NG[77 ] = (RAM_DEPTH > 32'h9A00) ? int_DB_DETECT_NG[77 ] : 1'b0;
    assign sel_DB_DETECT_NG[78 ] = (RAM_DEPTH > 32'h9C00) ? int_DB_DETECT_NG[78 ] : 1'b0;
    assign sel_DB_DETECT_NG[79 ] = (RAM_DEPTH > 32'h9E00) ? int_DB_DETECT_NG[79 ] : 1'b0;
    assign sel_DB_DETECT_NG[80 ] = (RAM_DEPTH > 32'hA000) ? int_DB_DETECT_NG[80 ] : 1'b0;
    assign sel_DB_DETECT_NG[81 ] = (RAM_DEPTH > 32'hA200) ? int_DB_DETECT_NG[81 ] : 1'b0;
    assign sel_DB_DETECT_NG[82 ] = (RAM_DEPTH > 32'hA400) ? int_DB_DETECT_NG[82 ] : 1'b0;
    assign sel_DB_DETECT_NG[83 ] = (RAM_DEPTH > 32'hA600) ? int_DB_DETECT_NG[83 ] : 1'b0;
    assign sel_DB_DETECT_NG[84 ] = (RAM_DEPTH > 32'hA800) ? int_DB_DETECT_NG[84 ] : 1'b0;
    assign sel_DB_DETECT_NG[85 ] = (RAM_DEPTH > 32'hAA00) ? int_DB_DETECT_NG[85 ] : 1'b0;
    assign sel_DB_DETECT_NG[86 ] = (RAM_DEPTH > 32'hAC00) ? int_DB_DETECT_NG[86 ] : 1'b0;
    assign sel_DB_DETECT_NG[87 ] = (RAM_DEPTH > 32'hAE00) ? int_DB_DETECT_NG[87 ] : 1'b0;
    assign sel_DB_DETECT_NG[88 ] = (RAM_DEPTH > 32'hB000) ? int_DB_DETECT_NG[88 ] : 1'b0;
    assign sel_DB_DETECT_NG[89 ] = (RAM_DEPTH > 32'hB200) ? int_DB_DETECT_NG[89 ] : 1'b0;
    assign sel_DB_DETECT_NG[90 ] = (RAM_DEPTH > 32'hB400) ? int_DB_DETECT_NG[90 ] : 1'b0;
    assign sel_DB_DETECT_NG[91 ] = (RAM_DEPTH > 32'hB600) ? int_DB_DETECT_NG[91 ] : 1'b0;
    assign sel_DB_DETECT_NG[92 ] = (RAM_DEPTH > 32'hB800) ? int_DB_DETECT_NG[92 ] : 1'b0;
    assign sel_DB_DETECT_NG[93 ] = (RAM_DEPTH > 32'hBA00) ? int_DB_DETECT_NG[93 ] : 1'b0;
    assign sel_DB_DETECT_NG[94 ] = (RAM_DEPTH > 32'hBC00) ? int_DB_DETECT_NG[94 ] : 1'b0;
    assign sel_DB_DETECT_NG[95 ] = (RAM_DEPTH > 32'hBE00) ? int_DB_DETECT_NG[95 ] : 1'b0;
    assign sel_DB_DETECT_NG[96 ] = (RAM_DEPTH > 32'hC000) ? int_DB_DETECT_NG[96 ] : 1'b0;
    assign sel_DB_DETECT_NG[97 ] = (RAM_DEPTH > 32'hC200) ? int_DB_DETECT_NG[97 ] : 1'b0;
    assign sel_DB_DETECT_NG[98 ] = (RAM_DEPTH > 32'hC400) ? int_DB_DETECT_NG[98 ] : 1'b0;
    assign sel_DB_DETECT_NG[99 ] = (RAM_DEPTH > 32'hC600) ? int_DB_DETECT_NG[99 ] : 1'b0;
    assign sel_DB_DETECT_NG[100] = (RAM_DEPTH > 32'hC800) ? int_DB_DETECT_NG[100] : 1'b0;
    assign sel_DB_DETECT_NG[101] = (RAM_DEPTH > 32'hCA00) ? int_DB_DETECT_NG[101] : 1'b0;
    assign sel_DB_DETECT_NG[102] = (RAM_DEPTH > 32'hCC00) ? int_DB_DETECT_NG[102] : 1'b0;
    assign sel_DB_DETECT_NG[103] = (RAM_DEPTH > 32'hCE00) ? int_DB_DETECT_NG[103] : 1'b0;
    assign sel_DB_DETECT_NG[104] = (RAM_DEPTH > 32'hD000) ? int_DB_DETECT_NG[104] : 1'b0;
    assign sel_DB_DETECT_NG[105] = (RAM_DEPTH > 32'hD200) ? int_DB_DETECT_NG[105] : 1'b0;
    assign sel_DB_DETECT_NG[106] = (RAM_DEPTH > 32'hD400) ? int_DB_DETECT_NG[106] : 1'b0;
    assign sel_DB_DETECT_NG[107] = (RAM_DEPTH > 32'hD600) ? int_DB_DETECT_NG[107] : 1'b0;
    assign sel_DB_DETECT_NG[108] = (RAM_DEPTH > 32'hD800) ? int_DB_DETECT_NG[108] : 1'b0;
    assign sel_DB_DETECT_NG[109] = (RAM_DEPTH > 32'hDA00) ? int_DB_DETECT_NG[109] : 1'b0;
    assign sel_DB_DETECT_NG[110] = (RAM_DEPTH > 32'hDC00) ? int_DB_DETECT_NG[110] : 1'b0;
    assign sel_DB_DETECT_NG[111] = (RAM_DEPTH > 32'hDE00) ? int_DB_DETECT_NG[111] : 1'b0;
    assign sel_DB_DETECT_NG[112] = (RAM_DEPTH > 32'hE000) ? int_DB_DETECT_NG[112] : 1'b0;
    assign sel_DB_DETECT_NG[113] = (RAM_DEPTH > 32'hE200) ? int_DB_DETECT_NG[113] : 1'b0;
    assign sel_DB_DETECT_NG[114] = (RAM_DEPTH > 32'hE400) ? int_DB_DETECT_NG[114] : 1'b0;
    assign sel_DB_DETECT_NG[115] = (RAM_DEPTH > 32'hE600) ? int_DB_DETECT_NG[115] : 1'b0;
    assign sel_DB_DETECT_NG[116] = (RAM_DEPTH > 32'hE800) ? int_DB_DETECT_NG[116] : 1'b0;
    assign sel_DB_DETECT_NG[117] = (RAM_DEPTH > 32'hEA00) ? int_DB_DETECT_NG[117] : 1'b0;
    assign sel_DB_DETECT_NG[118] = (RAM_DEPTH > 32'hEC00) ? int_DB_DETECT_NG[118] : 1'b0;
    assign sel_DB_DETECT_NG[119] = (RAM_DEPTH > 32'hEE00) ? int_DB_DETECT_NG[119] : 1'b0;
    assign sel_DB_DETECT_NG[120] = (RAM_DEPTH > 32'hF000) ? int_DB_DETECT_NG[120] : 1'b0;
    assign sel_DB_DETECT_NG[121] = (RAM_DEPTH > 32'hF200) ? int_DB_DETECT_NG[121] : 1'b0;
    assign sel_DB_DETECT_NG[122] = (RAM_DEPTH > 32'hF400) ? int_DB_DETECT_NG[122] : 1'b0;
    assign sel_DB_DETECT_NG[123] = (RAM_DEPTH > 32'hF600) ? int_DB_DETECT_NG[123] : 1'b0;
    assign sel_DB_DETECT_NG[124] = (RAM_DEPTH > 32'hF800) ? int_DB_DETECT_NG[124] : 1'b0;
    assign sel_DB_DETECT_NG[125] = (RAM_DEPTH > 32'hFA00) ? int_DB_DETECT_NG[125] : 1'b0;
    assign sel_DB_DETECT_NG[126] = (RAM_DEPTH > 32'hFC00) ? int_DB_DETECT_NG[126] : 1'b0;
    assign sel_DB_DETECT_NG[127] = (RAM_DEPTH > 32'hFE00) ? int_DB_DETECT_NG[127] : 1'b0;

    wire \SB_CORRECT[0] , \SB_CORRECT[1] , \SB_CORRECT[2] , 
        \SB_CORRECT[3] , \SB_CORRECT[4] , \SB_CORRECT[5] , 
        \SB_CORRECT[6] , \SB_CORRECT[7] , \SB_CORRECT[8] , 
        \SB_CORRECT[9] , \SB_CORRECT[10] , \SB_CORRECT[11] , 
        \SB_CORRECT[12] , \SB_CORRECT[13] , \SB_CORRECT[14] , 
        \SB_CORRECT[15] , \SB_CORRECT[16] , \SB_CORRECT[17] , 
        \SB_CORRECT[18] , \SB_CORRECT[19] , \SB_CORRECT[20] , 
        \SB_CORRECT[21] , \SB_CORRECT[22] , \SB_CORRECT[23] , 
        \SB_CORRECT[24] , \SB_CORRECT[25] , \SB_CORRECT[26] , 
        \SB_CORRECT[27] , \SB_CORRECT[28] , \SB_CORRECT[29] , 
        \SB_CORRECT[30] , \SB_CORRECT[31] , \SB_CORRECT[32] , 
        \SB_CORRECT[33] , \SB_CORRECT[34] , \SB_CORRECT[35] , 
        \SB_CORRECT[36] , \SB_CORRECT[37] , \SB_CORRECT[38] , 
        \SB_CORRECT[39] , \SB_CORRECT[40] , \SB_CORRECT[41] , 
        \SB_CORRECT[42] , \SB_CORRECT[43] , \SB_CORRECT[44] , 
        \SB_CORRECT[45] , \SB_CORRECT[46] , \SB_CORRECT[47] , 
        \SB_CORRECT[48] , \SB_CORRECT[49] , \SB_CORRECT[50] , 
        \SB_CORRECT[51] , \SB_CORRECT[52] , \SB_CORRECT[53] , 
        \SB_CORRECT[54] , \SB_CORRECT[55] , \SB_CORRECT[56] , 
        \SB_CORRECT[57] , \SB_CORRECT[58] , \SB_CORRECT[59] , 
        \SB_CORRECT[60] , \SB_CORRECT[61] , \SB_CORRECT[62] , 
        \SB_CORRECT[63] , \SB_CORRECT[64] , \SB_CORRECT[65] , 
        \SB_CORRECT[66] , \SB_CORRECT[67] , \SB_CORRECT[68] , 
        \SB_CORRECT[69] , \SB_CORRECT[70] , \SB_CORRECT[71] , 
        \SB_CORRECT[72] , \SB_CORRECT[73] , \SB_CORRECT[74] , 
        \SB_CORRECT[75] , \SB_CORRECT[76] , \SB_CORRECT[77] , 
        \SB_CORRECT[78] , \SB_CORRECT[79] , \SB_CORRECT[80] , 
        \SB_CORRECT[81] , \SB_CORRECT[82] , \SB_CORRECT[83] , 
        \SB_CORRECT[84] , \SB_CORRECT[85] , \SB_CORRECT[86] , 
        \SB_CORRECT[87] , \SB_CORRECT[88] , \SB_CORRECT[89] , 
        \SB_CORRECT[90] , \SB_CORRECT[91] , \SB_CORRECT[92] , 
        \SB_CORRECT[93] , \SB_CORRECT[94] , \SB_CORRECT[95] , 
        \SB_CORRECT[96] , \SB_CORRECT[97] , \SB_CORRECT[98] , 
        \SB_CORRECT[99] , \SB_CORRECT[100] , 
        \SB_CORRECT[101] , \SB_CORRECT[102] , 
        \SB_CORRECT[103] , \SB_CORRECT[104] , 
        \SB_CORRECT[105] , \SB_CORRECT[106] , 
        \SB_CORRECT[107] , \SB_CORRECT[108] , 
        \SB_CORRECT[109] , \SB_CORRECT[110] , 
        \SB_CORRECT[111] , \SB_CORRECT[112] , 
        \SB_CORRECT[113] , \SB_CORRECT[114] , 
        \SB_CORRECT[115] , \SB_CORRECT[116] , 
        \SB_CORRECT[117] , \SB_CORRECT[118] , 
        \SB_CORRECT[119] , \SB_CORRECT[120] , 
        \SB_CORRECT[121] , \SB_CORRECT[122] , 
        \SB_CORRECT[123] , \SB_CORRECT[124] , 
        \SB_CORRECT[125] , \SB_CORRECT[126] , 
        \SB_CORRECT[127] , \DB_DETECT[0] , \DB_DETECT[1] , 
        \DB_DETECT[2] , \DB_DETECT[3] , \DB_DETECT[4] , 
        \DB_DETECT[5] , \DB_DETECT[6] , \DB_DETECT[7] , 
        \DB_DETECT[8] , \DB_DETECT[9] , \DB_DETECT[10] , 
        \DB_DETECT[11] , \DB_DETECT[12] , \DB_DETECT[13] , 
        \DB_DETECT[14] , \DB_DETECT[15] , \DB_DETECT[16] , 
        \DB_DETECT[17] , \DB_DETECT[18] , \DB_DETECT[19] , 
        \DB_DETECT[20] , \DB_DETECT[21] , \DB_DETECT[22] , 
        \DB_DETECT[23] , \DB_DETECT[24] , \DB_DETECT[25] , 
        \DB_DETECT[26] , \DB_DETECT[27] , \DB_DETECT[28] , 
        \DB_DETECT[29] , \DB_DETECT[30] , \DB_DETECT[31] , 
        \DB_DETECT[32] , \DB_DETECT[33] , \DB_DETECT[34] , 
        \DB_DETECT[35] , \DB_DETECT[36] , \DB_DETECT[37] , 
        \DB_DETECT[38] , \DB_DETECT[39] , \DB_DETECT[40] , 
        \DB_DETECT[41] , \DB_DETECT[42] , \DB_DETECT[43] , 
        \DB_DETECT[44] , \DB_DETECT[45] , \DB_DETECT[46] , 
        \DB_DETECT[47] , \DB_DETECT[48] , \DB_DETECT[49] , 
        \DB_DETECT[50] , \DB_DETECT[51] , \DB_DETECT[52] , 
        \DB_DETECT[53] , \DB_DETECT[54] , \DB_DETECT[55] , 
        \DB_DETECT[56] , \DB_DETECT[57] , \DB_DETECT[58] , 
        \DB_DETECT[59] , \DB_DETECT[60] , \DB_DETECT[61] , 
        \DB_DETECT[62] , \DB_DETECT[63] , \DB_DETECT[64] , 
        \DB_DETECT[65] , \DB_DETECT[66] , \DB_DETECT[67] , 
        \DB_DETECT[68] , \DB_DETECT[69] , \DB_DETECT[70] , 
        \DB_DETECT[71] , \DB_DETECT[72] , \DB_DETECT[73] , 
        \DB_DETECT[74] , \DB_DETECT[75] , \DB_DETECT[76] , 
        \DB_DETECT[77] , \DB_DETECT[78] , \DB_DETECT[79] , 
        \DB_DETECT[80] , \DB_DETECT[81] , \DB_DETECT[82] , 
        \DB_DETECT[83] , \DB_DETECT[84] , \DB_DETECT[85] , 
        \DB_DETECT[86] , \DB_DETECT[87] , \DB_DETECT[88] , 
        \DB_DETECT[89] , \DB_DETECT[90] , \DB_DETECT[91] , 
        \DB_DETECT[92] , \DB_DETECT[93] , \DB_DETECT[94] , 
        \DB_DETECT[95] , \DB_DETECT[96] , \DB_DETECT[97] , 
        \DB_DETECT[98] , \DB_DETECT[99] , \DB_DETECT[100] , 
        \DB_DETECT[101] , \DB_DETECT[102] , \DB_DETECT[103] , 
        \DB_DETECT[104] , \DB_DETECT[105] , \DB_DETECT[106] , 
        \DB_DETECT[107] , \DB_DETECT[108] , \DB_DETECT[109] , 
        \DB_DETECT[110] , \DB_DETECT[111] , \DB_DETECT[112] , 
        \DB_DETECT[113] , \DB_DETECT[114] , \DB_DETECT[115] , 
        \DB_DETECT[116] , \DB_DETECT[117] , \DB_DETECT[118] , 
        \DB_DETECT[119] , \DB_DETECT[120] , \DB_DETECT[121] , 
        \DB_DETECT[122] , \DB_DETECT[123] , \DB_DETECT[124] , 
        \DB_DETECT[125] , \DB_DETECT[126] , \DB_DETECT[127] , 
        \BLKX0[0] , 
        \BLKY0[0] , \BLKY0_pipe[0] , \BLKY0_pipe[1] , \BLKX1[0] , 
        \BLKY1[0] , \BLKY1_pipe[0] , \BLKY1_pipe[1] , \BLKX2[0] , 
        \BLKX2[1] , \BLKX2[2] , \BLKX2[3] , \BLKX2[4] , \BLKX2[5] , 
        \BLKX2[6] , \BLKX2[7] , \BLKX2[8] , \BLKX2[9] , \BLKX2[10] , 
        \BLKX2[11] , \BLKX2[12] , \BLKX2[13] , \BLKX2[14] , 
        \BLKX2[15] , \BLKX2[16] , \BLKX2[17] , \BLKX2[18] , 
        \BLKX2[19] , \BLKX2[20] , \BLKX2[21] , \BLKX2[22] , 
        \BLKX2[23] , \BLKX2[24] , \BLKX2[25] , \BLKX2[26] , 
        \BLKX2[27] , \BLKX2[28] , \BLKX2[29] , \BLKX2[30] , 
        \BLKX2[31] , \BLKY2[0] , \BLKY2[1] , \BLKY2[2] , \BLKY2[3] , 
        \BLKY2[4] , \BLKY2[5] , \BLKY2[6] , \BLKY2[7] , \BLKY2[8] , 
        \BLKY2[9] , \BLKY2[10] , \BLKY2[11] , \BLKY2[12] , \BLKY2[13] , 
        \BLKY2[14] , \BLKY2[15] , \BLKY2[16] , \BLKY2[17] , 
        \BLKY2[18] , \BLKY2[19] , \BLKY2[20] , \BLKY2[21] , 
        \BLKY2[22] , \BLKY2[23] , \BLKY2[24] , \BLKY2[25] , 
        \BLKY2[26] , \BLKY2[27] , \BLKY2[28] , \BLKY2[29] , 
        \BLKY2[30] , \BLKY2[31] , \BLKY2_pipe[0] , \BLKY2_pipe[1] , 
        \BLKY2_pipe[2] , \BLKY2_pipe[3] , \BLKY2_pipe[4] , 
        \BLKY2_pipe[5] , \BLKY2_pipe[6] , \BLKY2_pipe[7] , 
        \BLKY2_pipe[8] , \BLKY2_pipe[9] , \BLKY2_pipe[10] , 
        \BLKY2_pipe[11] , \BLKY2_pipe[12] , \BLKY2_pipe[13] , 
        \BLKY2_pipe[14] , \BLKY2_pipe[15] , \BLKY2_pipe[16] , 
        \BLKY2_pipe[17] , \BLKY2_pipe[18] , \BLKY2_pipe[19] , 
        \BLKY2_pipe[20] , \BLKY2_pipe[21] , \BLKY2_pipe[22] , 
        \BLKY2_pipe[23] , \BLKY2_pipe[24] , \BLKY2_pipe[25] , 
        \BLKY2_pipe[26] , \BLKY2_pipe[27] , \BLKY2_pipe[28] , 
        \BLKY2_pipe[29] , \BLKY2_pipe[30] , \BLKY2_pipe[31] , 
        CFG3_16_Y, 
        CFG3_15_Y, CFG3_0_Y, CFG3_19_Y, CFG3_18_Y, CFG3_11_Y, CFG3_1_Y, 
        CFG3_21_Y, CFG3_2_Y, CFG3_20_Y, CFG3_9_Y, CFG3_3_Y, OR4_752_Y, 
        OR4_679_Y, OR4_946_Y, OR4_1046_Y, OR4_898_Y, OR4_427_Y, 
        OR4_906_Y, OR4_379_Y, OR4_922_Y, OR4_772_Y, OR4_1252_Y, 
        OR4_239_Y, OR4_1056_Y, OR4_1323_Y, OR4_843_Y, OR4_192_Y, 
        OR4_853_Y, OR4_1083_Y, OR4_1259_Y, OR4_716_Y, OR4_1181_Y, 
        OR4_171_Y, OR4_981_Y, OR4_1261_Y, OR4_770_Y, OR4_114_Y, 
        OR4_789_Y, OR4_1014_Y, OR4_1189_Y, OR4_976_Y, OR4_58_Y, 
        OR4_446_Y, OR4_1267_Y, OR4_122_Y, OR4_1048_Y, OR4_391_Y, 
        OR4_1060_Y, OR4_1290_Y, OR4_61_Y, OR4_1074_Y, OR4_143_Y, 
        OR2_15_Y, OR4_176_Y, OR4_831_Y, OR4_1203_Y, OR4_1327_Y, 
        OR4_298_Y, OR4_1052_Y, OR4_206_Y, OR4_852_Y, OR4_643_Y, 
        OR4_1250_Y, OR4_312_Y, OR4_1191_Y, OR4_4_Y, OR4_499_Y, 
        OR4_1168_Y, OR4_1389_Y, OR4_955_Y, OR4_734_Y, OR4_502_Y, 
        OR4_519_Y, OR4_967_Y, OR4_470_Y, OR4_665_Y, OR4_1165_Y, 
        OR4_456_Y, OR4_657_Y, OR4_246_Y, OR4_19_Y, OR4_1174_Y, 
        OR4_857_Y, OR4_1334_Y, OR4_805_Y, OR4_1024_Y, OR4_117_Y, 
        OR4_783_Y, OR4_1007_Y, OR4_587_Y, OR4_373_Y, OR4_123_Y, 
        OR4_987_Y, OR4_76_Y, OR2_23_Y, OR4_71_Y, OR4_378_Y, OR4_1003_Y, 
        OR4_482_Y, OR4_1350_Y, OR4_1041_Y, OR4_1363_Y, OR4_586_Y, 
        OR4_577_Y, OR4_429_Y, OR4_407_Y, OR4_125_Y, OR4_498_Y, 
        OR4_347_Y, OR4_1236_Y, OR4_285_Y, OR4_1253_Y, OR4_809_Y, 
        OR4_850_Y, OR4_730_Y, OR4_715_Y, OR4_457_Y, OR4_799_Y, 
        OR4_652_Y, OR4_142_Y, OR4_580_Y, OR4_170_Y, OR4_1130_Y, 
        OR4_1187_Y, OR4_1374_Y, OR4_1357_Y, OR4_1072_Y, OR4_55_Y, 
        OR4_1291_Y, OR4_767_Y, OR4_1234_Y, OR4_784_Y, OR4_375_Y, 
        OR4_425_Y, OR4_824_Y, OR4_804_Y, OR2_16_Y, OR4_331_Y, 
        OR4_710_Y, OR4_599_Y, OR4_706_Y, OR4_417_Y, OR4_856_Y, 
        OR4_1231_Y, OR4_467_Y, OR4_561_Y, OR4_359_Y, OR4_803_Y, 
        OR4_1205_Y, OR4_628_Y, OR4_886_Y, OR4_434_Y, OR4_1155_Y, 
        OR4_454_Y, OR4_655_Y, OR4_811_Y, OR4_740_Y, OR4_1207_Y, 
        OR4_197_Y, OR4_1012_Y, OR4_1283_Y, OR4_801_Y, OR4_148_Y, 
        OR4_817_Y, OR4_1040_Y, OR4_1219_Y, OR4_634_Y, OR4_1091_Y, 
        OR4_95_Y, OR4_905_Y, OR4_1180_Y, OR4_694_Y, OR4_48_Y, 
        OR4_717_Y, OR4_938_Y, OR4_1101_Y, OR4_735_Y, OR4_1204_Y, 
        OR2_5_Y, OR4_686_Y, OR4_845_Y, OR4_513_Y, OR4_1031_Y, 
        OR4_210_Y, OR4_297_Y, OR4_733_Y, OR4_284_Y, OR4_910_Y, 
        OR4_718_Y, OR4_1186_Y, OR4_173_Y, OR4_984_Y, OR4_1264_Y, 
        OR4_778_Y, OR4_116_Y, OR4_794_Y, OR4_1021_Y, OR4_1193_Y, 
        OR4_871_Y, OR4_1348_Y, OR4_339_Y, OR4_1162_Y, OR4_33_Y, 
        OR4_945_Y, OR4_300_Y, OR4_959_Y, OR4_1196_Y, OR4_1356_Y, 
        OR4_541_Y, OR4_989_Y, OR4_1388_Y, OR4_807_Y, OR4_1073_Y, 
        OR4_603_Y, OR4_1341_Y, OR4_620_Y, OR4_833_Y, OR4_996_Y, 
        OR4_1057_Y, OR4_121_Y, OR2_14_Y, OR4_525_Y, OR4_1286_Y, 
        OR4_134_Y, OR4_216_Y, OR4_1208_Y, OR4_773_Y, OR4_848_Y, 
        OR4_1111_Y, OR4_219_Y, OR4_207_Y, OR4_658_Y, OR4_146_Y, 
        OR4_358_Y, OR4_839_Y, OR4_120_Y, OR4_349_Y, OR4_1318_Y, 
        OR4_1093_Y, OR4_844_Y, OR4_948_Y, OR4_30_Y, OR4_892_Y, 
        OR4_1115_Y, OR4_217_Y, OR4_868_Y, OR4_1102_Y, OR4_673_Y, 
        OR4_466_Y, OR4_220_Y, OR4_1215_Y, OR4_282_Y, OR4_1149_Y, 
        OR4_1367_Y, OR4_465_Y, OR4_1126_Y, OR4_1358_Y, OR4_924_Y, 
        OR4_698_Y, OR4_471_Y, OR4_1278_Y, OR4_348_Y, OR2_29_Y, 
        OR4_325_Y, OR4_15_Y, OR4_1310_Y, OR4_1067_Y, OR4_867_Y, 
        OR4_1351_Y, OR4_552_Y, OR4_1120_Y, OR4_613_Y, OR4_1391_Y, 
        OR4_462_Y, OR4_1333_Y, OR4_149_Y, OR4_637_Y, OR4_1309_Y, 
        OR4_137_Y, OR4_1114_Y, OR4_877_Y, OR4_640_Y, OR4_1076_Y, 
        OR4_152_Y, OR4_1027_Y, OR4_1248_Y, OR4_340_Y, OR4_1004_Y, 
        OR4_1243_Y, OR4_797_Y, OR4_576_Y, OR4_343_Y, OR4_979_Y, 
        OR4_60_Y, OR4_926_Y, OR4_1138_Y, OR4_245_Y, OR4_907_Y, 
        OR4_1127_Y, OR4_707_Y, OR4_494_Y, OR4_249_Y, OR4_744_Y, 
        OR4_1220_Y, OR2_21_Y, OR4_223_Y, OR4_1319_Y, OR4_866_Y, 
        OR4_1146_Y, OR4_621_Y, OR4_1094_Y, OR4_978_Y, OR4_421_Y, 
        OR4_221_Y, OR4_263_Y, OR4_700_Y, OR4_1087_Y, OR4_523_Y, 
        OR4_774_Y, OR4_318_Y, OR4_1038_Y, OR4_336_Y, OR4_554_Y, 
        OR4_709_Y, OR4_1360_Y, OR4_422_Y, OR4_788_Y, OR4_236_Y, 
        OR4_500_Y, OR4_29_Y, OR4_749_Y, OR4_47_Y, OR4_269_Y, OR4_431_Y, 
        OR4_911_Y, OR4_1375_Y, OR4_365_Y, OR4_1194_Y, OR4_63_Y, 
        OR4_969_Y, OR4_316_Y, OR4_985_Y, OR4_1225_Y, OR4_1384_Y, 
        OR4_1185_Y, OR4_244_Y, OR2_19_Y, OR4_324_Y, OR4_261_Y, 
        OR4_283_Y, OR4_1245_Y, OR4_779_Y, OR4_1023_Y, OR4_1018_Y, 
        OR4_1260_Y, OR4_653_Y, OR4_670_Y, OR4_654_Y, OR4_390_Y, 
        OR4_747_Y, OR4_594_Y, OR4_99_Y, OR4_529_Y, OR4_106_Y, 
        OR4_1071_Y, OR4_1121_Y, OR4_601_Y, OR4_583_Y, OR4_320_Y, 
        OR4_672_Y, OR4_528_Y, OR4_16_Y, OR4_469_Y, OR4_43_Y, OR4_998_Y, 
        OR4_1045_Y, OR4_627_Y, OR4_607_Y, OR4_345_Y, OR4_695_Y, 
        OR4_556_Y, OR4_49_Y, OR4_491_Y, OR4_70_Y, OR4_1028_Y, 
        OR4_1068_Y, OR4_203_Y, OR4_182_Y, OR2_33_Y, OR4_873_Y, 
        OR4_834_Y, OR4_646_Y, OR4_31_Y, OR4_1136_Y, OR4_562_Y, 
        OR4_847_Y, OR4_162_Y, OR4_265_Y, OR4_559_Y, OR4_1015_Y, 
        OR4_509_Y, OR4_711_Y, OR4_1216_Y, OR4_492_Y, OR4_696_Y, 
        OR4_295_Y, OR4_69_Y, OR4_1222_Y, OR4_521_Y, OR4_971_Y, 
        OR4_472_Y, OR4_667_Y, OR4_1170_Y, OR4_458_Y, OR4_659_Y, 
        OR4_250_Y, OR4_22_Y, OR4_1176_Y, OR4_327_Y, OR4_771_Y, 
        OR4_278_Y, OR4_483_Y, OR4_960_Y, OR4_259_Y, OR4_476_Y, 
        OR4_56_Y, OR4_1228_Y, OR4_961_Y, OR4_1088_Y, OR4_164_Y, 
        OR2_25_Y, OR4_299_Y, OR4_951_Y, OR4_1311_Y, OR4_54_Y, 
        OR4_408_Y, OR4_1177_Y, OR4_321_Y, OR4_972_Y, OR4_756_Y, 
        OR4_781_Y, OR4_760_Y, OR4_50_Y, OR4_448_Y, OR4_691_Y, 
        OR4_900_Y, OR4_739_Y, OR4_442_Y, OR4_302_Y, OR4_403_Y, 
        OR4_80_Y, OR4_53_Y, OR4_708_Y, OR4_1112_Y, OR4_1377_Y, 
        OR4_188_Y, OR4_23_Y, OR4_1104_Y, OR4_953_Y, OR4_1062_Y, 
        OR4_433_Y, OR4_402_Y, OR4_1059_Y, OR4_78_Y, OR4_338_Y, 
        OR4_539_Y, OR4_377_Y, OR4_74_Y, OR4_1313_Y, OR4_35_Y, 
        OR4_550_Y, OR4_524_Y, OR2_28_Y, OR4_1086_Y, OR4_367_Y, 
        OR4_894_Y, OR4_510_Y, OR4_254_Y, OR4_1047_Y, OR4_1116_Y, 
        OR4_436_Y, OR4_1223_Y, OR4_757_Y, OR4_1239_Y, OR4_704_Y, 
        OR4_918_Y, OR4_20_Y, OR4_683_Y, OR4_902_Y, OR4_495_Y, 
        OR4_275_Y, OR4_24_Y, OR4_39_Y, OR4_504_Y, OR4_1379_Y, 
        OR4_194_Y, OR4_675_Y, OR4_1364_Y, OR4_184_Y, OR4_1157_Y, 
        OR4_927_Y, OR4_680_Y, OR4_571_Y, OR4_1035_Y, OR4_522_Y, 
        OR4_726_Y, OR4_1237_Y, OR4_507_Y, OR4_719_Y, OR4_310_Y, 
        OR4_91_Y, OR4_1240_Y, OR4_186_Y, OR4_639_Y, OR2_2_Y, OR4_800_Y, 
        OR4_1272_Y, OR4_869_Y, OR4_671_Y, OR4_1332_Y, OR4_202_Y, 
        OR4_1008_Y, OR4_846_Y, OR4_374_Y, OR4_829_Y, OR4_1297_Y, 
        OR4_301_Y, OR4_1118_Y, OR4_1383_Y, OR4_896_Y, OR4_248_Y, 
        OR4_920_Y, OR4_1140_Y, OR4_1301_Y, OR4_1296_Y, OR4_360_Y, 
        OR4_741_Y, OR4_178_Y, OR4_451_Y, OR4_1368_Y, OR4_689_Y, 
        OR4_1386_Y, OR4_212_Y, OR4_371_Y, OR4_914_Y, OR4_1376_Y, 
        OR4_366_Y, OR4_1195_Y, OR4_66_Y, OR4_970_Y, OR4_317_Y, 
        OR4_986_Y, OR4_1227_Y, OR4_1385_Y, OR4_705_Y, OR4_1173_Y, 
        OR2_4_Y, OR4_518_Y, OR4_1263_Y, OR4_765_Y, OR4_256_Y, 
        OR4_1361_Y, OR4_865_Y, OR4_59_Y, OR4_650_Y, OR4_1080_Y, 
        OR4_937_Y, OR4_656_Y, OR4_1070_Y, OR4_745_Y, OR4_798_Y, 
        OR4_526_Y, OR4_585_Y, OR4_994_Y, OR4_880_Y, OR4_816_Y, 
        OR4_296_Y, OR4_12_Y, OR4_432_Y, OR4_102_Y, OR4_155_Y, 
        OR4_1275_Y, OR4_1336_Y, OR4_355_Y, OR4_240_Y, OR4_174_Y, 
        OR4_1202_Y, OR4_917_Y, OR4_1335_Y, OR4_1002_Y, OR4_1058_Y, 
        OR4_775_Y, OR4_842_Y, OR4_1268_Y, OR4_1147_Y, OR4_1075_Y, 
        OR4_663_Y, OR4_394_Y, OR2_22_Y, OR4_642_Y, OR4_9_Y, OR4_266_Y, 
        OR4_329_Y, OR4_1315_Y, OR4_893_Y, OR4_963_Y, OR4_1235_Y, 
        OR4_335_Y, OR4_1148_Y, OR4_1123_Y, OR4_399_Y, OR4_780_Y, 
        OR4_1053_Y, OR4_1269_Y, OR4_1098_Y, OR4_776_Y, OR4_645_Y, 
        OR4_750_Y, OR4_512_Y, OR4_490_Y, OR4_1151_Y, OR4_153_Y, 
        OR4_428_Y, OR4_622_Y, OR4_468_Y, OR4_151_Y, OR4_11_Y, 
        OR4_112_Y, OR4_753_Y, OR4_728_Y, OR4_8_Y, OR4_404_Y, OR4_661_Y, 
        OR4_858_Y, OR4_702_Y, OR4_398_Y, OR4_267_Y, OR4_369_Y, 
        OR4_819_Y, OR4_792_Y, OR2_0_Y, OR4_447_Y, OR4_129_Y, OR4_37_Y, 
        OR4_1197_Y, OR4_988_Y, OR4_77_Y, OR4_660_Y, OR4_1246_Y, 
        OR4_731_Y, OR4_936_Y, OR4_915_Y, OR4_190_Y, OR4_574_Y, 
        OR4_840_Y, OR4_1051_Y, OR4_882_Y, OR4_573_Y, OR4_450_Y, 
        OR4_546_Y, OR4_631_Y, OR4_605_Y, OR4_1280_Y, OR4_292_Y, 
        OR4_545_Y, OR4_748_Y, OR4_579_Y, OR4_289_Y, OR4_132_Y, 
        OR4_247_Y, OR4_538_Y, OR4_515_Y, OR4_1190_Y, OR4_187_Y, 
        OR4_460_Y, OR4_648_Y, OR4_497_Y, OR4_179_Y, OR4_41_Y, 
        OR4_144_Y, OR4_309_Y, OR4_287_Y, OR2_24_Y, CFG3_13_Y, CFG3_8_Y, 
        CFG3_14_Y, CFG3_5_Y, CFG3_6_Y, CFG3_22_Y, CFG3_10_Y, CFG3_23_Y, 
        CFG3_12_Y, CFG3_4_Y, CFG3_17_Y, CFG3_7_Y, OR4_1122_Y, 
        OR4_1299_Y, OR4_912_Y, OR4_724_Y, OR4_1276_Y, OR4_17_Y, 
        OR4_118_Y, OR4_26_Y, OR4_814_Y, OR4_1153_Y, OR4_222_Y, 
        OR4_595_Y, OR4_36_Y, OR4_308_Y, OR4_1232_Y, OR4_557_Y, 
        OR4_1247_Y, OR4_72_Y, OR4_227_Y, OR4_1330_Y, OR4_396_Y, 
        OR4_768_Y, OR4_214_Y, OR4_478_Y, OR4_5_Y, OR4_725_Y, OR4_18_Y, 
        OR4_241_Y, OR4_400_Y, OR4_940_Y, OR4_10_Y, OR4_397_Y, 
        OR4_1230_Y, OR4_96_Y, OR4_1005_Y, OR4_351_Y, OR4_1025_Y, 
        OR4_1258_Y, OR4_14_Y, OR4_755_Y, OR4_1226_Y, OR2_7_Y, 
        OR4_992_Y, OR4_954_Y, OR4_758_Y, OR4_140_Y, OR4_1262_Y, 
        OR4_677_Y, OR4_962_Y, OR4_286_Y, OR4_372_Y, OR4_108_Y, 
        OR4_97_Y, OR4_751_Y, OR4_1150_Y, OR4_25_Y, OR4_230_Y, OR4_75_Y, 
        OR4_1143_Y, OR4_993_Y, OR4_1117_Y, OR4_84_Y, OR4_57_Y, 
        OR4_712_Y, OR4_1113_Y, OR4_1381_Y, OR4_191_Y, OR4_27_Y, 
        OR4_1110_Y, OR4_956_Y, OR4_1065_Y, OR4_1274_Y, OR4_1254_Y, 
        OR4_520_Y, OR4_908_Y, OR4_1188_Y, OR4_1390_Y, OR4_1233_Y, 
        OR4_901_Y, OR4_761_Y, OR4_859_Y, OR4_644_Y, OR4_611_Y, 
        OR2_31_Y, OR4_1218_Y, OR4_485_Y, OR4_1011_Y, OR4_618_Y, 
        OR4_364_Y, OR4_1171_Y, OR4_1241_Y, OR4_543_Y, OR4_1331_Y, 
        OR4_319_Y, OR4_304_Y, OR4_952_Y, OR4_1362_Y, OR4_229_Y, 
        OR4_444_Y, OR4_279_Y, OR4_1359_Y, OR4_1221_Y, OR4_1314_Y, 
        OR4_973_Y, OR4_949_Y, OR4_234_Y, OR4_623_Y, OR4_883_Y, 
        OR4_1095_Y, OR4_933_Y, OR4_614_Y, OR4_487_Y, OR4_581_Y, 
        OR4_124_Y, OR4_104_Y, OR4_764_Y, OR4_1169_Y, OR4_45_Y, 
        OR4_251_Y, OR4_92_Y, OR4_1164_Y, OR4_1016_Y, OR4_1125_Y, 
        OR4_1124_Y, OR4_1105_Y, OR2_9_Y, OR4_1211_Y, OR4_713_Y, 
        OR4_7_Y, OR4_602_Y, OR4_966_Y, OR4_1277_Y, OR4_34_Y, 
        OR4_1042_Y, OR4_1082_Y, OR4_861_Y, OR4_1340_Y, OR4_812_Y, 
        OR4_1029_Y, OR4_126_Y, OR4_790_Y, OR4_1017_Y, OR4_593_Y, 
        OR4_382_Y, OR4_130_Y, OR4_393_Y, OR4_841_Y, OR4_337_Y, 
        OR4_542_Y, OR4_1034_Y, OR4_314_Y, OR4_531_Y, OR4_110_Y, 
        OR4_1287_Y, OR4_1037_Y, OR4_1063_Y, OR4_135_Y, OR4_1006_Y, 
        OR4_1238_Y, OR4_326_Y, OR4_983_Y, OR4_1224_Y, OR4_782_Y, 
        OR4_564_Y, OR4_332_Y, OR4_293_Y, OR4_738_Y, OR2_8_Y, OR4_181_Y, 
        OR4_449_Y, OR4_787_Y, OR4_1061_Y, OR4_441_Y, OR4_1229_Y, 
        OR4_759_Y, OR4_305_Y, OR4_714_Y, OR4_218_Y, OR4_662_Y, 
        OR4_1050_Y, OR4_493_Y, OR4_743_Y, OR4_290_Y, OR4_999_Y, 
        OR4_306_Y, OR4_516_Y, OR4_666_Y, OR4_475_Y, OR4_921_Y, 
        OR4_1308_Y, OR4_737_Y, OR4_995_Y, OR4_532_Y, OR4_1270_Y, 
        OR4_551_Y, OR4_763_Y, OR4_925_Y, OR4_820_Y, OR4_1289_Y, 
        OR4_291_Y, OR4_1107_Y, OR4_1373_Y, OR4_889_Y, OR4_237_Y, 
        OR4_909_Y, OR4_1128_Y, OR4_1294_Y, OR4_1099_Y, OR4_169_Y, 
        OR2_17_Y, OR4_1142_Y, OR4_1305_Y, OR4_854_Y, OR4_1129_Y, 
        OR4_1090_Y, OR4_1079_Y, OR4_990_Y, OR4_1345_Y, OR4_209_Y, 
        OR4_1183_Y, OR4_242_Y, OR4_619_Y, OR4_65_Y, OR4_322_Y, 
        OR4_1251_Y, OR4_572_Y, OR4_1266_Y, OR4_94_Y, OR4_253_Y, 
        OR4_1342_Y, OR4_409_Y, OR4_777_Y, OR4_225_Y, OR4_489_Y, 
        OR4_13_Y, OR4_736_Y, OR4_32_Y, OR4_260_Y, OR4_416_Y, OR4_891_Y, 
        OR4_1366_Y, OR4_354_Y, OR4_1182_Y, OR4_52_Y, OR4_958_Y, 
        OR4_311_Y, OR4_975_Y, OR4_1213_Y, OR4_1370_Y, OR4_1167_Y, 
        OR4_231_Y, OR2_18_Y, OR4_1010_Y, OR4_1338_Y, OR4_567_Y, 
        OR4_44_Y, OR4_899_Y, OR4_606_Y, OR4_919_Y, OR4_163_Y, 
        OR4_150_Y, OR4_687_Y, OR4_1154_Y, OR4_633_Y, OR4_836_Y, 
        OR4_1344_Y, OR4_608_Y, OR4_827_Y, OR4_424_Y, OR4_196_Y, 
        OR4_1349_Y, OR4_1001_Y, OR4_88_Y, OR4_943_Y, OR4_1163_Y, 
        OR4_270_Y, OR4_932_Y, OR4_1152_Y, OR4_727_Y, OR4_511_Y, 
        OR4_273_Y, OR4_257_Y, OR4_701_Y, OR4_193_Y, OR4_406_Y, 
        OR4_885_Y, OR4_175_Y, OR4_395_Y, OR4_1369_Y, OR4_1137_Y, 
        OR4_890_Y, OR4_1109_Y, OR4_177_Y, OR2_26_Y, OR4_723_Y, 
        OR4_368_Y, OR4_313_Y, OR4_277_Y, OR4_1198_Y, OR4_904_Y, 
        OR4_881_Y, OR4_356_Y, OR4_111_Y, OR4_410_Y, OR4_851_Y, 
        OR4_350_Y, OR4_558_Y, OR4_1044_Y, OR4_334_Y, OR4_548_Y, 
        OR4_119_Y, OR4_1298_Y, OR4_1049_Y, OR4_40_Y, OR4_505_Y, 
        OR4_1380_Y, OR4_195_Y, OR4_676_Y, OR4_1365_Y, OR4_185_Y, 
        OR4_1158_Y, OR4_928_Y, OR4_681_Y, OR4_1387_Y, OR4_459_Y, 
        OR4_1328_Y, OR4_139_Y, OR4_630_Y, OR4_1302_Y, OR4_127_Y, 
        OR4_1106_Y, OR4_863_Y, OR4_632_Y, OR4_1337_Y, OR4_405_Y, 
        OR2_30_Y, OR4_1316_Y, OR4_822_Y, OR4_113_Y, OR4_720_Y, 
        OR4_1089_Y, OR4_1393_Y, OR4_145_Y, OR4_1166_Y, OR4_1212_Y, 
        OR4_437_Y, OR4_411_Y, OR4_1064_Y, OR4_83_Y, OR4_341_Y, 
        OR4_544_Y, OR4_384_Y, OR4_79_Y, OR4_1321_Y, OR4_38_Y, 
        OR4_1339_Y, OR4_1307_Y, OR4_575_Y, OR4_968_Y, OR4_1255_Y, 
        OR4_67_Y, OR4_1288_Y, OR4_964_Y, OR4_825_Y, OR4_939_Y, 
        OR4_615_Y, OR4_588_Y, OR4_1271_Y, OR4_276_Y, OR4_530_Y, 
        OR4_732_Y, OR4_568_Y, OR4_271_Y, OR4_115_Y, OR4_232_Y, 
        OR4_1242_Y, OR4_1209_Y, OR2_13_Y, OR4_1214_Y, OR4_1013_Y, 
        OR4_385_Y, OR4_569_Y, OR4_769_Y, OR4_496_Y, OR4_268_Y, 
        OR4_328_Y, OR4_294_Y, OR4_862_Y, OR4_1343_Y, OR4_813_Y, 
        OR4_1030_Y, OR4_128_Y, OR4_791_Y, OR4_1019_Y, OR4_596_Y, 
        OR4_383_Y, OR4_133_Y, OR4_688_Y, OR4_1156_Y, OR4_635_Y, 
        OR4_837_Y, OR4_1346_Y, OR4_609_Y, OR4_828_Y, OR4_426_Y, 
        OR4_198_Y, OR4_1352_Y, OR4_62_Y, OR4_517_Y, OR4_1_Y, OR4_215_Y, 
        OR4_690_Y, OR4_1378_Y, OR4_204_Y, OR4_1178_Y, OR4_941_Y, 
        OR4_697_Y, OR4_258_Y, OR4_703_Y, OR2_6_Y, OR4_323_Y, OR4_977_Y, 
        OR4_51_Y, OR4_243_Y, OR4_189_Y, OR4_636_Y, OR4_333_Y, 
        OR4_330_Y, OR4_280_Y, OR4_353_Y, OR4_796_Y, OR4_1199_Y, 
        OR4_617_Y, OR4_872_Y, OR4_423_Y, OR4_1145_Y, OR4_443_Y, 
        OR4_647_Y, OR4_802_Y, OR4_1009_Y, OR4_93_Y, OR4_473_Y, 
        OR4_1293_Y, OR4_165_Y, OR4_1077_Y, OR4_430_Y, OR4_1100_Y, 
        OR4_1322_Y, OR4_98_Y, OR4_86_Y, OR4_527_Y, OR4_916_Y, 
        OR4_352_Y, OR4_604_Y, OR4_138_Y, OR4_855_Y, OR4_159_Y, 
        OR4_380_Y, OR4_535_Y, OR4_281_Y, OR4_721_Y, OR2_27_Y, 
        OR4_1279_Y, OR4_1217_Y, OR4_1244_Y, OR4_785_Y, OR4_357_Y, 
        OR4_584_Y, OR4_578_Y, OR4_806_Y, OR4_228_Y, OR4_942_Y, 
        OR4_21_Y, OR4_887_Y, OR4_1108_Y, OR4_211_Y, OR4_860_Y, 
        OR4_1092_Y, OR4_668_Y, OR4_461_Y, OR4_213_Y, OR4_864_Y, 
        OR4_1347_Y, OR4_815_Y, OR4_1032_Y, OR4_131_Y, OR4_795_Y, 
        OR4_1022_Y, OR4_597_Y, OR4_386_Y, OR4_136_Y, OR4_895_Y, 
        OR4_1371_Y, OR4_838_Y, OR4_1054_Y, OR4_161_Y, OR4_818_Y, 
        OR4_1043_Y, OR4_625_Y, OR4_412_Y, OR4_167_Y, OR4_481_Y, 
        OR4_930_Y, OR2_11_Y, OR4_1131_Y, OR4_64_Y, OR4_682_Y, 
        OR4_154_Y, OR4_1020_Y, OR4_722_Y, OR4_1033_Y, OR4_288_Y, 
        OR4_274_Y, OR4_252_Y, OR4_224_Y, OR4_876_Y, OR4_1284_Y, 
        OR4_157_Y, OR4_361_Y, OR4_200_Y, OR4_1281_Y, OR4_1133_Y, 
        OR4_1256_Y, OR4_560_Y, OR4_533_Y, OR4_1210_Y, OR4_208_Y, 
        OR4_477_Y, OR4_669_Y, OR4_514_Y, OR4_205_Y, OR4_68_Y, 
        OR4_172_Y, OR4_1200_Y, OR4_1172_Y, OR4_455_Y, OR4_826_Y, 
        OR4_1103_Y, OR4_1304_Y, OR4_1141_Y, OR4_823_Y, OR4_685_Y, 
        OR4_786_Y, OR4_651_Y, OR4_629_Y, OR2_32_Y, OR4_1055_Y, 
        OR4_272_Y, OR4_453_Y, OR4_591_Y, OR4_160_Y, OR4_418_Y, 
        OR4_168_Y, OR4_875_Y, OR4_105_Y, OR4_1085_Y, OR4_156_Y, 
        OR4_540_Y, OR4_1372_Y, OR4_238_Y, OR4_1160_Y, OR4_501_Y, 
        OR4_1179_Y, OR4_3_Y, OR4_166_Y, OR4_307_Y, OR4_746_Y, 
        OR4_1134_Y, OR4_563_Y, OR4_821_Y, OR4_362_Y, OR4_1084_Y, 
        OR4_381_Y, OR4_590_Y, OR4_754_Y, OR4_480_Y, OR4_923_Y, 
        OR4_1312_Y, OR4_742_Y, OR4_1000_Y, OR4_536_Y, OR4_1273_Y, 
        OR4_555_Y, OR4_766_Y, OR4_935_Y, OR4_626_Y, OR4_1081_Y, 
        OR2_1_Y, OR4_832_Y, OR4_486_Y, OR4_435_Y, OR4_388_Y, 
        OR4_1303_Y, OR4_1026_Y, OR4_997_Y, OR4_474_Y, OR4_233_Y, 
        OR4_1355_Y, OR4_1326_Y, OR4_589_Y, OR4_982_Y, OR4_1265_Y, 
        OR4_82_Y, OR4_1300_Y, OR4_980_Y, OR4_835_Y, OR4_947_Y, 
        OR4_974_Y, OR4_950_Y, OR4_235_Y, OR4_624_Y, OR4_884_Y, 
        OR4_1096_Y, OR4_934_Y, OR4_616_Y, OR4_488_Y, OR4_582_Y, 
        OR4_931_Y, OR4_897_Y, OR4_183_Y, OR4_570_Y, OR4_830_Y, 
        OR4_1039_Y, OR4_870_Y, OR4_565_Y, OR4_438_Y, OR4_537_Y, 
        OR4_874_Y, OR4_849_Y, OR2_3_Y, OR4_1392_Y, OR4_109_Y, 
        OR4_592_Y, OR4_1249_Y, OR4_729_Y, OR4_1192_Y, OR4_303_Y, 
        OR4_100_Y, OR4_315_Y, OR4_762_Y, OR4_957_Y, OR4_553_Y, 
        OR4_1036_Y, OR4_534_Y, OR4_1206_Y, OR4_678_Y, OR4_1184_Y, 
        OR4_692_Y, OR4_90_Y, OR4_879_Y, OR4_1078_Y, OR4_664_Y, 
        OR4_1159_Y, OR4_649_Y, OR4_1317_Y, OR4_793_Y, OR4_1295_Y, 
        OR4_810_Y, OR4_199_Y, OR4_1382_Y, OR4_180_Y, OR4_1161_Y, 
        OR4_264_Y, OR4_1139_Y, OR4_420_Y, OR4_1292_Y, OR4_392_Y, 
        OR4_1306_Y, OR4_674_Y, OR4_612_Y, OR4_808_Y, OR2_10_Y, 
        OR4_1320_Y, OR4_1132_Y, OR4_503_Y, OR4_684_Y, OR4_888_Y, 
        OR4_598_Y, OR4_376_Y, OR4_452_Y, OR4_401_Y, OR4_439_Y, 
        OR4_413_Y, OR4_1066_Y, OR4_87_Y, OR4_344_Y, OR4_547_Y, 
        OR4_387_Y, OR4_81_Y, OR4_1324_Y, OR4_42_Y, OR4_255_Y, 
        OR4_226_Y, OR4_878_Y, OR4_1285_Y, OR4_158_Y, OR4_363_Y, 
        OR4_201_Y, OR4_1282_Y, OR4_1135_Y, OR4_1257_Y, OR4_991_Y, 
        OR4_965_Y, OR4_262_Y, OR4_641_Y, OR4_903_Y, OR4_1119_Y, 
        OR4_944_Y, OR4_638_Y, OR4_506_Y, OR4_600_Y, OR4_1201_Y, 
        OR4_1175_Y, OR2_12_Y, OR4_2_Y, OR4_1325_Y, OR4_1353_Y, 
        OR4_913_Y, OR4_479_Y, OR4_699_Y, OR4_693_Y, OR4_929_Y, 
        OR4_342_Y, OR4_508_Y, OR4_484_Y, OR4_1144_Y, OR4_147_Y, 
        OR4_419_Y, OR4_610_Y, OR4_463_Y, OR4_141_Y, OR4_6_Y, OR4_107_Y, 
        OR4_445_Y, OR4_415_Y, OR4_1069_Y, OR4_89_Y, OR4_346_Y, 
        OR4_549_Y, OR4_389_Y, OR4_85_Y, OR4_1329_Y, OR4_46_Y, 
        OR4_464_Y, OR4_440_Y, OR4_1097_Y, OR4_103_Y, OR4_370_Y, 
        OR4_566_Y, OR4_414_Y, OR4_101_Y, OR4_1354_Y, OR4_73_Y, 
        OR4_28_Y, OR4_0_Y, OR2_20_Y, ADLIB_GND, VCC, GND, ADLIB_VCC;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign ADLIB_GND = GND_power_net1;
    assign GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign ADLIB_VCC = VCC_power_net1;
    
    OR4 OR4_700 (.A(sel_R_DATA_TEMPR88[5] ), .B(sel_R_DATA_TEMPR89[5] ), .C(sel_R_DATA_TEMPR90[5] ), .D(sel_R_DATA_TEMPR91[5] ), .Y(OR4_700_Y));
    OR4 OR4_399 (.A(sel_R_DATA_TEMPR92[16] ), .B(sel_R_DATA_TEMPR93[16] ), 
        .C(sel_R_DATA_TEMPR94[16] ), .D(sel_R_DATA_TEMPR95[16] ), .Y(
        OR4_399_Y));
    OR4 OR4_1188 (.A(sel_R_DATA_TEMPR52[12] ), .B(sel_R_DATA_TEMPR53[12] ), 
        .C(sel_R_DATA_TEMPR54[12] ), .D(sel_R_DATA_TEMPR55[12] ), .Y(
        OR4_1188_Y));
    OR4 OR4_420 (.A(\DB_DETECT[56] ), .B(\DB_DETECT[57] ), .C(
        \DB_DETECT[58] ), .D(\DB_DETECT[59] ), .Y(OR4_420_Y));
    OR4 OR4_738 (.A(sel_R_DATA_TEMPR80[24] ), .B(sel_R_DATA_TEMPR81[24] ), 
        .C(sel_R_DATA_TEMPR82[24] ), .D(sel_R_DATA_TEMPR83[24] ), .Y(
        OR4_738_Y));
    OR4 OR4_1141 (.A(sel_R_DATA_TEMPR60[10] ), .B(sel_R_DATA_TEMPR61[10] ), 
        .C(sel_R_DATA_TEMPR62[10] ), .D(sel_R_DATA_TEMPR63[10] ), .Y(
        OR4_1141_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[1]  (.A(CFG3_15_Y), .B(CFG3_2_Y)
        , .Y(\BLKY2[1] ));
    OR4 OR4_402 (.A(sel_R_DATA_TEMPR40[17] ), .B(sel_R_DATA_TEMPR41[17] ), 
        .C(sel_R_DATA_TEMPR42[17] ), .D(sel_R_DATA_TEMPR43[17] ), .Y(
        OR4_402_Y));
    AND4 \AND4DB_DETECT[117]  (.A(sel_DB_DETECT_NG[117] ), .B(
        \BLKY2_pipe[29] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[117] ));
    OR4 OR4_384 (.A(sel_R_DATA_TEMPR108[14] ), .B(sel_R_DATA_TEMPR109[14] ), 
        .C(sel_R_DATA_TEMPR110[14] ), .D(sel_R_DATA_TEMPR111[14] ), .Y(
        OR4_384_Y));
    OR4 OR4_373 (.A(sel_R_DATA_TEMPR68[27] ), .B(sel_R_DATA_TEMPR69[27] ), 
        .C(sel_R_DATA_TEMPR70[27] ), .D(sel_R_DATA_TEMPR71[27] ), .Y(
        OR4_373_Y));
    OR4 OR4_770 (.A(sel_R_DATA_TEMPR16[2] ), .B(sel_R_DATA_TEMPR17[2] ), .C(sel_R_DATA_TEMPR18[2] ), .D(sel_R_DATA_TEMPR19[2] ), .Y(OR4_770_Y));
    OR4 OR4_253 (.A(sel_R_DATA_TEMPR120[0] ), .B(sel_R_DATA_TEMPR121[0] ), 
        .C(sel_R_DATA_TEMPR122[0] ), .D(sel_R_DATA_TEMPR123[0] ), .Y(
        OR4_253_Y));
    OR4 OR4_1331 (.A(OR4_1164_Y), .B(OR4_1016_Y), .C(OR4_1125_Y), .D(
        OR4_1124_Y), .Y(OR4_1331_Y));
    OR4 OR4_1253 (.A(sel_R_DATA_TEMPR112[30] ), .B(sel_R_DATA_TEMPR113[30] ), 
        .C(sel_R_DATA_TEMPR114[30] ), .D(sel_R_DATA_TEMPR115[30] ), .Y(
        OR4_1253_Y));
    OR4 OR4_409 (.A(sel_R_DATA_TEMPR0[0] ), .B(sel_R_DATA_TEMPR1[0] ), .C(sel_R_DATA_TEMPR2[0] ), .D(sel_R_DATA_TEMPR3[0] ), .Y(OR4_409_Y));
    OR4 OR4_472 (.A(sel_R_DATA_TEMPR4[22] ), .B(sel_R_DATA_TEMPR5[22] ), .C(sel_R_DATA_TEMPR6[22] ), .D(sel_R_DATA_TEMPR7[22] ), .Y(OR4_472_Y));
    OR4 OR4_181 (.A(OR4_441_Y), .B(OR4_1229_Y), .C(OR4_759_Y), .D(
        OR4_305_Y), .Y(OR4_181_Y));
    OR4 OR4_961 (.A(sel_R_DATA_TEMPR72[22] ), .B(sel_R_DATA_TEMPR73[22] ), 
        .C(sel_R_DATA_TEMPR74[22] ), .D(sel_R_DATA_TEMPR75[22] ), .Y(
        OR4_961_Y));
    OR4 OR4_106 (.A(sel_R_DATA_TEMPR112[31] ), .B(sel_R_DATA_TEMPR113[31] ), 
        .C(sel_R_DATA_TEMPR114[31] ), .D(sel_R_DATA_TEMPR115[31] ), .Y(
        OR4_106_Y));
    AND4 \AND4DB_DETECT[30]  (.A(sel_DB_DETECT_NG[30] ), .B(
        \BLKY2_pipe[7] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[30] ));
    AND4 \AND4DB_DETECT[14]  (.A(sel_DB_DETECT_NG[14] ), .B(
        \BLKY2_pipe[3] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[14] ));
    OR4 OR4_958 (.A(sel_R_DATA_TEMPR56[0] ), .B(sel_R_DATA_TEMPR57[0] ), .C(sel_R_DATA_TEMPR58[0] ), .D(sel_R_DATA_TEMPR59[0] ), .Y(OR4_958_Y));
    OR4 OR4_83 (.A(sel_R_DATA_TEMPR96[14] ), .B(sel_R_DATA_TEMPR97[14] ), .C(sel_R_DATA_TEMPR98[14] ), .D(sel_R_DATA_TEMPR99[14] ), .Y(OR4_83_Y));
    OR4 OR4_479 (.A(OR4_415_Y), .B(OR4_1069_Y), .C(OR4_89_Y), .D(
        OR4_346_Y), .Y(OR4_479_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[22]  (.A(CFG3_10_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[22] ));
    OR4 OR4_837 (.A(sel_R_DATA_TEMPR8[28] ), .B(sel_R_DATA_TEMPR9[28] ), .C(sel_R_DATA_TEMPR10[28] ), .D(sel_R_DATA_TEMPR11[28] ), .Y(OR4_837_Y));
    OR4 OR4_138 (.A(sel_R_DATA_TEMPR56[6] ), .B(sel_R_DATA_TEMPR57[6] ), .C(sel_R_DATA_TEMPR58[6] ), .D(sel_R_DATA_TEMPR59[6] ), .Y(OR4_138_Y));
    OR4 OR4_934 (.A(sel_R_DATA_TEMPR20[13] ), .B(sel_R_DATA_TEMPR21[13] ), 
        .C(sel_R_DATA_TEMPR22[13] ), .D(sel_R_DATA_TEMPR23[13] ), .Y(
        OR4_934_Y));
    OR4 OR4_176 (.A(OR4_298_Y), .B(OR4_1052_Y), .C(OR4_206_Y), .D(
        OR4_852_Y), .Y(OR4_176_Y));
    OR4 OR4_610 (.A(sel_R_DATA_TEMPR104[11] ), .B(sel_R_DATA_TEMPR105[11] ), 
        .C(sel_R_DATA_TEMPR106[11] ), .D(sel_R_DATA_TEMPR107[11] ), .Y(
        OR4_610_Y));
    OR4 OR4_481 (.A(sel_R_DATA_TEMPR76[21] ), .B(sel_R_DATA_TEMPR77[21] ), 
        .C(sel_R_DATA_TEMPR78[21] ), .D(sel_R_DATA_TEMPR79[21] ), .Y(
        OR4_481_Y));
    OR4 OR4_1216 (.A(sel_R_DATA_TEMPR100[22] ), .B(sel_R_DATA_TEMPR101[22] ), 
        .C(sel_R_DATA_TEMPR102[22] ), .D(sel_R_DATA_TEMPR103[22] ), .Y(
        OR4_1216_Y));
    AND4 \AND4SB_CORRECT[108]  (.A(sel_SB_CORRECT_NG[108] ), .B(
        \BLKY2_pipe[27] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[108] ));
    AND4 \AND4SB_CORRECT[70]  (.A(sel_SB_CORRECT_NG[70] ), .B(
        \BLKY2_pipe[17] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[70] ));
    OR4 OR4_488 (.A(sel_R_DATA_TEMPR28[13] ), .B(sel_R_DATA_TEMPR29[13] ), 
        .C(sel_R_DATA_TEMPR30[13] ), .D(sel_R_DATA_TEMPR31[13] ), .Y(
        OR4_488_Y));
    OR4 OR4_1072 (.A(sel_R_DATA_TEMPR44[30] ), .B(sel_R_DATA_TEMPR45[30] ), 
        .C(sel_R_DATA_TEMPR46[30] ), .D(sel_R_DATA_TEMPR47[30] ), .Y(
        OR4_1072_Y));
    OR4 OR4_308 (.A(sel_R_DATA_TEMPR100[1] ), .B(sel_R_DATA_TEMPR101[1] ), 
        .C(sel_R_DATA_TEMPR102[1] ), .D(sel_R_DATA_TEMPR103[1] ), .Y(
        OR4_308_Y));
    OR4 OR4_1159 (.A(\DB_DETECT[8] ), .B(\DB_DETECT[9] ), .C(
        \DB_DETECT[10] ), .D(\DB_DETECT[11] ), .Y(OR4_1159_Y));
    OR4 OR4_317 (.A(sel_R_DATA_TEMPR60[7] ), .B(sel_R_DATA_TEMPR61[7] ), .C(sel_R_DATA_TEMPR62[7] ), .D(sel_R_DATA_TEMPR63[7] ), .Y(OR4_317_Y));
    OR4 OR4_110 (.A(sel_R_DATA_TEMPR24[24] ), .B(sel_R_DATA_TEMPR25[24] ), 
        .C(sel_R_DATA_TEMPR26[24] ), .D(sel_R_DATA_TEMPR27[24] ), .Y(
        OR4_110_Y));
    OR4 OR4_848 (.A(OR4_220_Y), .B(OR4_1215_Y), .C(OR4_282_Y), .D(
        OR4_1149_Y), .Y(OR4_848_Y));
    OR4 OR4_1318 (.A(sel_R_DATA_TEMPR112[26] ), .B(sel_R_DATA_TEMPR113[26] ), 
        .C(sel_R_DATA_TEMPR114[26] ), .D(sel_R_DATA_TEMPR115[26] ), .Y(
        OR4_1318_Y));
    CFG3 #( .INIT(8'h1) )  CFG3_16 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_16_Y));
    OR4 OR4_1026 (.A(OR4_1096_Y), .B(OR4_934_Y), .C(OR4_616_Y), .D(
        OR4_488_Y), .Y(OR4_1026_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[8]  (.D(\BLKY2[8] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[8] ));
    OR4 OR4_658 (.A(sel_R_DATA_TEMPR88[26] ), .B(sel_R_DATA_TEMPR89[26] ), 
        .C(sel_R_DATA_TEMPR90[26] ), .D(sel_R_DATA_TEMPR91[26] ), .Y(
        OR4_658_Y));
    OR4 OR4_1045 (.A(sel_R_DATA_TEMPR32[31] ), .B(sel_R_DATA_TEMPR33[31] ), 
        .C(sel_R_DATA_TEMPR34[31] ), .D(sel_R_DATA_TEMPR35[31] ), .Y(
        OR4_1045_Y));
    OR4 OR4_799 (.A(sel_R_DATA_TEMPR8[30] ), .B(sel_R_DATA_TEMPR9[30] ), .C(sel_R_DATA_TEMPR10[30] ), .D(sel_R_DATA_TEMPR11[30] ), .Y(OR4_799_Y));
    OR4 OR4_378 (.A(OR4_577_Y), .B(OR4_429_Y), .C(OR4_407_Y), .D(
        OR4_125_Y), .Y(OR4_378_Y));
    OR4 OR4_2 (.A(OR4_479_Y), .B(OR4_699_Y), .C(OR4_693_Y), .D(
        OR4_929_Y), .Y(OR4_2_Y));
    OR4 OR4_718 (.A(OR4_121_Y), .B(OR2_14_Y), .C(sel_R_DATA_TEMPR86[8] ), 
        .D(sel_R_DATA_TEMPR87[8] ), .Y(OR4_718_Y));
    AND4 \AND4SB_CORRECT[29]  (.A(sel_SB_CORRECT_NG[29] ), .B(
        \BLKY2_pipe[7] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[29] ));
    OR4 OR4_329 (.A(OR4_776_Y), .B(OR4_645_Y), .C(OR4_750_Y), .D(
        OR4_512_Y), .Y(OR4_329_Y));
    AND4 \AND4SB_CORRECT[91]  (.A(sel_SB_CORRECT_NG[91] ), .B(
        \BLKY2_pipe[22] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[91] ));
    OR4 \OR4_R_DATA[29]  (.A(OR4_325_Y), .B(OR4_15_Y), .C(OR4_1310_Y), 
        .D(OR4_1067_Y), .Y(R_DATA[29]));
    OR4 OR4_894 (.A(OR4_918_Y), .B(OR4_20_Y), .C(OR4_683_Y), .D(
        OR4_902_Y), .Y(OR4_894_Y));
    OR4 OR4_765 (.A(OR4_745_Y), .B(OR4_798_Y), .C(OR4_526_Y), .D(
        OR4_585_Y), .Y(OR4_765_Y));
    OR4 OR4_667 (.A(sel_R_DATA_TEMPR8[22] ), .B(sel_R_DATA_TEMPR9[22] ), .C(sel_R_DATA_TEMPR10[22] ), .D(sel_R_DATA_TEMPR11[22] ), .Y(OR4_667_Y));
    OR4 OR4_652 (.A(sel_R_DATA_TEMPR12[30] ), .B(sel_R_DATA_TEMPR13[30] ), 
        .C(sel_R_DATA_TEMPR14[30] ), .D(sel_R_DATA_TEMPR15[30] ), .Y(
        OR4_652_Y));
    OR4 OR4_1321 (.A(sel_R_DATA_TEMPR116[14] ), .B(sel_R_DATA_TEMPR117[14] ), 
        .C(sel_R_DATA_TEMPR118[14] ), .D(sel_R_DATA_TEMPR119[14] ), .Y(
        OR4_1321_Y));
    OR4 OR4_766 (.A(sel_R_DATA_TEMPR68[4] ), .B(sel_R_DATA_TEMPR69[4] ), .C(sel_R_DATA_TEMPR70[4] ), .D(sel_R_DATA_TEMPR71[4] ), .Y(OR4_766_Y));
    OR4 OR4_593 (.A(sel_R_DATA_TEMPR112[24] ), .B(sel_R_DATA_TEMPR113[24] ), 
        .C(sel_R_DATA_TEMPR114[24] ), .D(sel_R_DATA_TEMPR115[24] ), .Y(
        OR4_593_Y));
    OR4 OR4_48 (.A(sel_R_DATA_TEMPR60[3] ), .B(sel_R_DATA_TEMPR61[3] ), .C(sel_R_DATA_TEMPR62[3] ), .D(sel_R_DATA_TEMPR63[3] ), .Y(OR4_48_Y));
    OR4 OR4_589 (.A(sel_R_DATA_TEMPR92[13] ), .B(sel_R_DATA_TEMPR93[13] ), 
        .C(sel_R_DATA_TEMPR94[13] ), .D(sel_R_DATA_TEMPR95[13] ), .Y(
        OR4_589_Y));
    OR2 OR2_33 (.A(sel_R_DATA_TEMPR84[31] ), .B(sel_R_DATA_TEMPR85[31] ), .Y(
        OR2_33_Y));
    OR4 OR4_109 (.A(OR4_315_Y), .B(OR4_762_Y), .C(OR4_957_Y), .D(
        OR4_553_Y), .Y(OR4_109_Y));
    OR2 OR2_15 (.A(sel_R_DATA_TEMPR84[2] ), .B(sel_R_DATA_TEMPR85[2] ), .Y(
        OR2_15_Y));
    AND4 \AND4SB_CORRECT[42]  (.A(sel_SB_CORRECT_NG[42] ), .B(
        \BLKY2_pipe[10] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[42] ));
    OR4 OR4_241 (.A(sel_R_DATA_TEMPR28[1] ), .B(sel_R_DATA_TEMPR29[1] ), .C(sel_R_DATA_TEMPR30[1] ), .D(sel_R_DATA_TEMPR31[1] ), .Y(OR4_241_Y));
    OR4 OR4_580 (.A(sel_R_DATA_TEMPR20[30] ), .B(sel_R_DATA_TEMPR21[30] ), 
        .C(sel_R_DATA_TEMPR22[30] ), .D(sel_R_DATA_TEMPR23[30] ), .Y(
        OR4_580_Y));
    AND4 \AND4SB_CORRECT[88]  (.A(sel_SB_CORRECT_NG[88] ), .B(
        \BLKY2_pipe[22] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[88] ));
    OR4 OR4_81 (.A(sel_R_DATA_TEMPR112[18] ), .B(sel_R_DATA_TEMPR113[18] ), 
        .C(sel_R_DATA_TEMPR114[18] ), .D(sel_R_DATA_TEMPR115[18] ), .Y(
        OR4_81_Y));
    OR4 OR4_1019 (.A(sel_R_DATA_TEMPR108[28] ), .B(sel_R_DATA_TEMPR109[28] ), 
        .C(sel_R_DATA_TEMPR110[28] ), .D(sel_R_DATA_TEMPR111[28] ), .Y(
        OR4_1019_Y));
    OR4 OR4_817 (.A(sel_R_DATA_TEMPR24[3] ), .B(sel_R_DATA_TEMPR25[3] ), .C(sel_R_DATA_TEMPR26[3] ), .D(sel_R_DATA_TEMPR27[3] ), .Y(OR4_817_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%94%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R94C0 (.A_DOUT({
        nc0, nc1, nc2, nc3, nc4,int_R_DATA_TEMPR94[31] , 
       int_R_DATA_TEMPR94[30] ,int_R_DATA_TEMPR94[29] , 
       int_R_DATA_TEMPR94[28] ,int_R_DATA_TEMPR94[27] , 
       int_R_DATA_TEMPR94[26] ,int_R_DATA_TEMPR94[25] , 
       int_R_DATA_TEMPR94[24] ,int_R_DATA_TEMPR94[23] , 
       int_R_DATA_TEMPR94[22] ,int_R_DATA_TEMPR94[21] , 
       int_R_DATA_TEMPR94[20] ,int_R_DATA_TEMPR94[19] , 
       int_R_DATA_TEMPR94[18] ,int_R_DATA_TEMPR94[17] }), .B_DOUT({nc5, 
        nc6, nc7,int_R_DATA_TEMPR94[16] ,int_R_DATA_TEMPR94[15] , 
       int_R_DATA_TEMPR94[14] ,int_R_DATA_TEMPR94[13] , 
       int_R_DATA_TEMPR94[12] ,int_R_DATA_TEMPR94[11] , 
       int_R_DATA_TEMPR94[10] ,int_R_DATA_TEMPR94[9] ,int_R_DATA_TEMPR94[8] , 
       int_R_DATA_TEMPR94[7] ,int_R_DATA_TEMPR94[6] ,int_R_DATA_TEMPR94[5] , 
       int_R_DATA_TEMPR94[4] ,int_R_DATA_TEMPR94[3] ,int_R_DATA_TEMPR94[2] , 
       int_R_DATA_TEMPR94[1] ,int_R_DATA_TEMPR94[0] }), .DB_DETECT( int_DB_DETECT_NG[94] ), .SB_CORRECT(int_SB_CORRECT_NG[94] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[94] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[23] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[23] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_118 (.A(OR4_400_Y), .B(OR4_940_Y), .C(OR4_10_Y), .D(
        OR4_397_Y), .Y(OR4_118_Y));
    OR4 OR4_914 (.A(sel_R_DATA_TEMPR36[7] ), .B(sel_R_DATA_TEMPR37[7] ), .C(sel_R_DATA_TEMPR38[7] ), .D(sel_R_DATA_TEMPR39[7] ), .Y(OR4_914_Y));
    OR4 \OR4_R_DATA[7]  (.A(OR4_800_Y), .B(OR4_1272_Y), .C(OR4_869_Y), 
        .D(OR4_671_Y), .Y(R_DATA[7]));
    AND4 \AND4DB_DETECT[12]  (.A(sel_DB_DETECT_NG[12] ), .B(
        \BLKY2_pipe[3] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[12] ));
    OR4 OR4_179 (.A(sel_R_DATA_TEMPR64[19] ), .B(sel_R_DATA_TEMPR65[19] ), 
        .C(sel_R_DATA_TEMPR66[19] ), .D(sel_R_DATA_TEMPR67[19] ), .Y(
        OR4_179_Y));
    OR4 OR4_1163 (.A(sel_R_DATA_TEMPR8[20] ), .B(sel_R_DATA_TEMPR9[20] ), .C(sel_R_DATA_TEMPR10[20] ), .D(sel_R_DATA_TEMPR11[20] ), .Y(OR4_1163_Y)
        );
    OR4 OR4_1156 (.A(sel_R_DATA_TEMPR0[28] ), .B(sel_R_DATA_TEMPR1[28] ), .C(sel_R_DATA_TEMPR2[28] ), .D(sel_R_DATA_TEMPR3[28] ), .Y(OR4_1156_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%8%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R8C0 (.A_DOUT({nc8, 
        nc9, nc10, nc11, nc12,int_R_DATA_TEMPR8[31] , 
       int_R_DATA_TEMPR8[30] ,int_R_DATA_TEMPR8[29] ,int_R_DATA_TEMPR8[28] , 
       int_R_DATA_TEMPR8[27] ,int_R_DATA_TEMPR8[26] ,int_R_DATA_TEMPR8[25] , 
       int_R_DATA_TEMPR8[24] ,int_R_DATA_TEMPR8[23] ,int_R_DATA_TEMPR8[22] , 
       int_R_DATA_TEMPR8[21] ,int_R_DATA_TEMPR8[20] ,int_R_DATA_TEMPR8[19] , 
       int_R_DATA_TEMPR8[18] ,int_R_DATA_TEMPR8[17] }), .B_DOUT({nc13, 
        nc14, nc15,int_R_DATA_TEMPR8[16] ,int_R_DATA_TEMPR8[15] , 
       int_R_DATA_TEMPR8[14] ,int_R_DATA_TEMPR8[13] ,int_R_DATA_TEMPR8[12] , 
       int_R_DATA_TEMPR8[11] ,int_R_DATA_TEMPR8[10] ,int_R_DATA_TEMPR8[9] , 
       int_R_DATA_TEMPR8[8] ,int_R_DATA_TEMPR8[7] ,int_R_DATA_TEMPR8[6] , 
       int_R_DATA_TEMPR8[5] ,int_R_DATA_TEMPR8[4] ,int_R_DATA_TEMPR8[3] , 
       int_R_DATA_TEMPR8[2] ,int_R_DATA_TEMPR8[1] ,int_R_DATA_TEMPR8[0] }), 
        .DB_DETECT(int_DB_DETECT_NG[8] ), .SB_CORRECT( int_SB_CORRECT_NG[8] ), .ACCESS_BUSY(\ACCESS_BUSY[8] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1251 (.A(sel_R_DATA_TEMPR104[0] ), .B(sel_R_DATA_TEMPR105[0] ), 
        .C(sel_R_DATA_TEMPR106[0] ), .D(sel_R_DATA_TEMPR107[0] ), .Y(
        OR4_1251_Y));
    OR4 OR4_901 (.A(sel_R_DATA_TEMPR64[12] ), .B(sel_R_DATA_TEMPR65[12] ), 
        .C(sel_R_DATA_TEMPR66[12] ), .D(sel_R_DATA_TEMPR67[12] ), .Y(
        OR4_901_Y));
    OR4 OR4_1158 (.A(sel_R_DATA_TEMPR24[23] ), .B(sel_R_DATA_TEMPR25[23] ), 
        .C(sel_R_DATA_TEMPR26[23] ), .D(sel_R_DATA_TEMPR27[23] ), .Y(
        OR4_1158_Y));
    AND4 \AND4SB_CORRECT[50]  (.A(sel_SB_CORRECT_NG[50] ), .B(
        \BLKY2_pipe[12] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[50] ));
    OR4 OR4_542 (.A(sel_R_DATA_TEMPR8[24] ), .B(sel_R_DATA_TEMPR9[24] ), .C(sel_R_DATA_TEMPR10[24] ), .D(sel_R_DATA_TEMPR11[24] ), .Y(OR4_542_Y));
    OR4 OR4_1132 (.A(OR4_401_Y), .B(OR4_439_Y), .C(OR4_413_Y), .D(
        OR4_1066_Y), .Y(OR4_1132_Y));
    OR4 OR4_855 (.A(sel_R_DATA_TEMPR60[6] ), .B(sel_R_DATA_TEMPR61[6] ), .C(sel_R_DATA_TEMPR62[6] ), .D(sel_R_DATA_TEMPR63[6] ), .Y(OR4_855_Y));
    AND4 \AND4SB_CORRECT[69]  (.A(sel_SB_CORRECT_NG[69] ), .B(
        \BLKY2_pipe[17] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[69] ));
    OR4 OR4_971 (.A(sel_R_DATA_TEMPR0[22] ), .B(sel_R_DATA_TEMPR1[22] ), .C(sel_R_DATA_TEMPR2[22] ), .D(sel_R_DATA_TEMPR3[22] ), .Y(OR4_971_Y));
    AND4 \AND4DB_DETECT[24]  (.A(sel_DB_DETECT_NG[24] ), .B(
        \BLKY2_pipe[6] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[24] ));
    OR4 OR4_729 (.A(OR4_1078_Y), .B(OR4_664_Y), .C(OR4_1159_Y), .D(
        OR4_649_Y), .Y(OR4_729_Y));
    OR4 \OR4_R_DATA[4]  (.A(OR4_1055_Y), .B(OR4_272_Y), .C(OR4_453_Y), 
        .D(OR4_591_Y), .Y(R_DATA[4]));
    OR4 OR4_135 (.A(sel_R_DATA_TEMPR40[24] ), .B(sel_R_DATA_TEMPR41[24] ), 
        .C(sel_R_DATA_TEMPR42[24] ), .D(sel_R_DATA_TEMPR43[24] ), .Y(
        OR4_135_Y));
    OR4 OR4_824 (.A(sel_R_DATA_TEMPR76[30] ), .B(sel_R_DATA_TEMPR77[30] ), 
        .C(sel_R_DATA_TEMPR78[30] ), .D(sel_R_DATA_TEMPR79[30] ), .Y(
        OR4_824_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[9]  (.A(CFG3_15_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[9] ));
    OR4 OR4_383 (.A(sel_R_DATA_TEMPR116[28] ), .B(sel_R_DATA_TEMPR117[28] ), 
        .C(sel_R_DATA_TEMPR118[28] ), .D(sel_R_DATA_TEMPR119[28] ), .Y(
        OR4_383_Y));
    OR4 OR4_1305 (.A(OR4_209_Y), .B(OR4_1183_Y), .C(OR4_242_Y), .D(
        OR4_619_Y), .Y(OR4_1305_Y));
    OR4 OR4_1140 (.A(sel_R_DATA_TEMPR116[7] ), .B(sel_R_DATA_TEMPR117[7] ), 
        .C(sel_R_DATA_TEMPR118[7] ), .D(sel_R_DATA_TEMPR119[7] ), .Y(
        OR4_1140_Y));
    OR4 OR4_780 (.A(sel_R_DATA_TEMPR96[16] ), .B(sel_R_DATA_TEMPR97[16] ), 
        .C(sel_R_DATA_TEMPR98[16] ), .D(sel_R_DATA_TEMPR99[16] ), .Y(
        OR4_780_Y));
    OR4 OR4_544 (.A(sel_R_DATA_TEMPR104[14] ), .B(sel_R_DATA_TEMPR105[14] ), 
        .C(sel_R_DATA_TEMPR106[14] ), .D(sel_R_DATA_TEMPR107[14] ), .Y(
        OR4_544_Y));
    OR2 OR2_31 (.A(sel_R_DATA_TEMPR84[12] ), .B(sel_R_DATA_TEMPR85[12] ), .Y(
        OR2_31_Y));
    OR4 OR4_267 (.A(sel_R_DATA_TEMPR68[16] ), .B(sel_R_DATA_TEMPR69[16] ), 
        .C(sel_R_DATA_TEMPR70[16] ), .D(sel_R_DATA_TEMPR71[16] ), .Y(
        OR4_267_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_9 (.A(R_EN), .B(R_ADDR[15]), .C(
        R_ADDR[14]), .Y(CFG3_9_Y));
    OR4 OR4_523 (.A(sel_R_DATA_TEMPR96[5] ), .B(sel_R_DATA_TEMPR97[5] ), .C(sel_R_DATA_TEMPR98[5] ), .D(sel_R_DATA_TEMPR99[5] ), .Y(OR4_523_Y));
    OR4 OR4_437 (.A(OR4_1209_Y), .B(OR2_13_Y), .C(sel_R_DATA_TEMPR86[14] )
        , .D(sel_R_DATA_TEMPR87[14] ), .Y(OR4_437_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%49%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R49C0 (.A_DOUT({
        nc16, nc17, nc18, nc19, nc20,int_R_DATA_TEMPR49[31] , 
       int_R_DATA_TEMPR49[30] ,int_R_DATA_TEMPR49[29] , 
       int_R_DATA_TEMPR49[28] ,int_R_DATA_TEMPR49[27] , 
       int_R_DATA_TEMPR49[26] ,int_R_DATA_TEMPR49[25] , 
       int_R_DATA_TEMPR49[24] ,int_R_DATA_TEMPR49[23] , 
       int_R_DATA_TEMPR49[22] ,int_R_DATA_TEMPR49[21] , 
       int_R_DATA_TEMPR49[20] ,int_R_DATA_TEMPR49[19] , 
       int_R_DATA_TEMPR49[18] ,int_R_DATA_TEMPR49[17] }), .B_DOUT({nc21, 
        nc22, nc23,int_R_DATA_TEMPR49[16] ,int_R_DATA_TEMPR49[15] , 
       int_R_DATA_TEMPR49[14] ,int_R_DATA_TEMPR49[13] , 
       int_R_DATA_TEMPR49[12] ,int_R_DATA_TEMPR49[11] , 
       int_R_DATA_TEMPR49[10] ,int_R_DATA_TEMPR49[9] ,int_R_DATA_TEMPR49[8] , 
       int_R_DATA_TEMPR49[7] ,int_R_DATA_TEMPR49[6] ,int_R_DATA_TEMPR49[5] , 
       int_R_DATA_TEMPR49[4] ,int_R_DATA_TEMPR49[3] ,int_R_DATA_TEMPR49[2] , 
       int_R_DATA_TEMPR49[1] ,int_R_DATA_TEMPR49[0] }), .DB_DETECT( int_DB_DETECT_NG[49] ), .SB_CORRECT(int_SB_CORRECT_NG[49] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[49] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[12] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4DB_DETECT[57]  (.A(sel_DB_DETECT_NG[57] ), .B(
        \BLKY2_pipe[14] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[57] ));
    OR4 OR4_942 (.A(OR4_930_Y), .B(OR2_11_Y), .C(sel_R_DATA_TEMPR86[21] ), 
        .D(sel_R_DATA_TEMPR87[21] ), .Y(OR4_942_Y));
    OR4 OR4_482 (.A(OR4_1253_Y), .B(OR4_809_Y), .C(OR4_850_Y), .D(
        OR4_730_Y), .Y(OR4_482_Y));
    OR4 OR4_167 (.A(sel_R_DATA_TEMPR72[21] ), .B(sel_R_DATA_TEMPR73[21] ), 
        .C(sel_R_DATA_TEMPR74[21] ), .D(sel_R_DATA_TEMPR75[21] ), .Y(
        OR4_167_Y));
    OR4 OR4_1193 (.A(sel_R_DATA_TEMPR120[8] ), .B(sel_R_DATA_TEMPR121[8] ), 
        .C(sel_R_DATA_TEMPR122[8] ), .D(sel_R_DATA_TEMPR123[8] ), .Y(
        OR4_1193_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%122%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R122C0 (.A_DOUT({
        nc24, nc25, nc26, nc27, nc28,int_R_DATA_TEMPR122[31] , 
       int_R_DATA_TEMPR122[30] ,int_R_DATA_TEMPR122[29] , 
       int_R_DATA_TEMPR122[28] ,int_R_DATA_TEMPR122[27] , 
       int_R_DATA_TEMPR122[26] ,int_R_DATA_TEMPR122[25] , 
       int_R_DATA_TEMPR122[24] ,int_R_DATA_TEMPR122[23] , 
       int_R_DATA_TEMPR122[22] ,int_R_DATA_TEMPR122[21] , 
       int_R_DATA_TEMPR122[20] ,int_R_DATA_TEMPR122[19] , 
       int_R_DATA_TEMPR122[18] ,int_R_DATA_TEMPR122[17] }), .B_DOUT({nc29, 
        nc30, nc31,int_R_DATA_TEMPR122[16] ,int_R_DATA_TEMPR122[15] , 
       int_R_DATA_TEMPR122[14] ,int_R_DATA_TEMPR122[13] , 
       int_R_DATA_TEMPR122[12] ,int_R_DATA_TEMPR122[11] , 
       int_R_DATA_TEMPR122[10] ,int_R_DATA_TEMPR122[9] , 
       int_R_DATA_TEMPR122[8] ,int_R_DATA_TEMPR122[7] , 
       int_R_DATA_TEMPR122[6] ,int_R_DATA_TEMPR122[5] , 
       int_R_DATA_TEMPR122[4] ,int_R_DATA_TEMPR122[3] , 
       int_R_DATA_TEMPR122[2] ,int_R_DATA_TEMPR122[1] , 
       int_R_DATA_TEMPR122[0] }), .DB_DETECT(int_DB_DETECT_NG[122] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[122] ), .ACCESS_BUSY(
        ACCESS_BUSY[122] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[30] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[30] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_705 (.A(sel_R_DATA_TEMPR76[7] ), .B(sel_R_DATA_TEMPR77[7] ), .C(sel_R_DATA_TEMPR78[7] ), .D(sel_R_DATA_TEMPR79[7] ), .Y(OR4_705_Y));
    OR4 OR4_607 (.A(sel_R_DATA_TEMPR40[31] ), .B(sel_R_DATA_TEMPR41[31] ), 
        .C(sel_R_DATA_TEMPR42[31] ), .D(sel_R_DATA_TEMPR43[31] ), .Y(
        OR4_607_Y));
    OR4 OR4_489 (.A(sel_R_DATA_TEMPR12[0] ), .B(sel_R_DATA_TEMPR13[0] ), .C(sel_R_DATA_TEMPR14[0] ), .D(sel_R_DATA_TEMPR15[0] ), .Y(OR4_489_Y));
    OR4 OR4_706 (.A(OR4_454_Y), .B(OR4_655_Y), .C(OR4_811_Y), .D(
        OR4_740_Y), .Y(OR4_706_Y));
    OR4 OR4_186 (.A(sel_R_DATA_TEMPR76[25] ), .B(sel_R_DATA_TEMPR77[25] ), 
        .C(sel_R_DATA_TEMPR78[25] ), .D(sel_R_DATA_TEMPR79[25] ), .Y(
        OR4_186_Y));
    OR4 OR4_775 (.A(\SB_CORRECT[56] ), .B(\SB_CORRECT[57] ), .C(
        \SB_CORRECT[58] ), .D(\SB_CORRECT[59] ), .Y(OR4_775_Y));
    OR4 OR4_677 (.A(OR4_191_Y), .B(OR4_27_Y), .C(OR4_1110_Y), .D(
        OR4_956_Y), .Y(OR4_677_Y));
    OR4 OR4_235 (.A(sel_R_DATA_TEMPR4[13] ), .B(sel_R_DATA_TEMPR5[13] ), .C(sel_R_DATA_TEMPR6[13] ), .D(sel_R_DATA_TEMPR7[13] ), .Y(OR4_235_Y));
    AND4 \AND4DB_DETECT[38]  (.A(sel_DB_DETECT_NG[38] ), .B(
        \BLKY2_pipe[9] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[38] ));
    OR4 OR4_341 (.A(sel_R_DATA_TEMPR100[14] ), .B(sel_R_DATA_TEMPR101[14] ), 
        .C(sel_R_DATA_TEMPR102[14] ), .D(sel_R_DATA_TEMPR103[14] ), .Y(
        OR4_341_Y));
    OR4 OR4_776 (.A(sel_R_DATA_TEMPR112[16] ), .B(sel_R_DATA_TEMPR113[16] ), 
        .C(sel_R_DATA_TEMPR114[16] ), .D(sel_R_DATA_TEMPR115[16] ), .Y(
        OR4_776_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[25]  (.D(\BLKY2[25] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[25] ));
    OR4 OR4_1122 (.A(OR4_1276_Y), .B(OR4_17_Y), .C(OR4_118_Y), .D(
        OR4_26_Y), .Y(OR4_1122_Y));
    OR4 OR4_763 (.A(sel_R_DATA_TEMPR28[9] ), .B(sel_R_DATA_TEMPR29[9] ), .C(sel_R_DATA_TEMPR30[9] ), .D(sel_R_DATA_TEMPR31[9] ), .Y(OR4_763_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%120%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R120C0 (.A_DOUT({
        nc32, nc33, nc34, nc35, nc36,int_R_DATA_TEMPR120[31] , 
       int_R_DATA_TEMPR120[30] ,int_R_DATA_TEMPR120[29] , 
       int_R_DATA_TEMPR120[28] ,int_R_DATA_TEMPR120[27] , 
       int_R_DATA_TEMPR120[26] ,int_R_DATA_TEMPR120[25] , 
       int_R_DATA_TEMPR120[24] ,int_R_DATA_TEMPR120[23] , 
       int_R_DATA_TEMPR120[22] ,int_R_DATA_TEMPR120[21] , 
       int_R_DATA_TEMPR120[20] ,int_R_DATA_TEMPR120[19] , 
       int_R_DATA_TEMPR120[18] ,int_R_DATA_TEMPR120[17] }), .B_DOUT({nc37, 
        nc38, nc39,int_R_DATA_TEMPR120[16] ,int_R_DATA_TEMPR120[15] , 
       int_R_DATA_TEMPR120[14] ,int_R_DATA_TEMPR120[13] , 
       int_R_DATA_TEMPR120[12] ,int_R_DATA_TEMPR120[11] , 
       int_R_DATA_TEMPR120[10] ,int_R_DATA_TEMPR120[9] , 
       int_R_DATA_TEMPR120[8] ,int_R_DATA_TEMPR120[7] , 
       int_R_DATA_TEMPR120[6] ,int_R_DATA_TEMPR120[5] , 
       int_R_DATA_TEMPR120[4] ,int_R_DATA_TEMPR120[3] , 
       int_R_DATA_TEMPR120[2] ,int_R_DATA_TEMPR120[1] , 
       int_R_DATA_TEMPR120[0] }), .DB_DETECT(int_DB_DETECT_NG[120] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[120] ), .ACCESS_BUSY(
        ACCESS_BUSY[120] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[30] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[30] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%123%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R123C0 (.A_DOUT({
        nc40, nc41, nc42, nc43, nc44,int_R_DATA_TEMPR123[31] , 
       int_R_DATA_TEMPR123[30] ,int_R_DATA_TEMPR123[29] , 
       int_R_DATA_TEMPR123[28] ,int_R_DATA_TEMPR123[27] , 
       int_R_DATA_TEMPR123[26] ,int_R_DATA_TEMPR123[25] , 
       int_R_DATA_TEMPR123[24] ,int_R_DATA_TEMPR123[23] , 
       int_R_DATA_TEMPR123[22] ,int_R_DATA_TEMPR123[21] , 
       int_R_DATA_TEMPR123[20] ,int_R_DATA_TEMPR123[19] , 
       int_R_DATA_TEMPR123[18] ,int_R_DATA_TEMPR123[17] }), .B_DOUT({nc45, 
        nc46, nc47,int_R_DATA_TEMPR123[16] ,int_R_DATA_TEMPR123[15] , 
       int_R_DATA_TEMPR123[14] ,int_R_DATA_TEMPR123[13] , 
       int_R_DATA_TEMPR123[12] ,int_R_DATA_TEMPR123[11] , 
       int_R_DATA_TEMPR123[10] ,int_R_DATA_TEMPR123[9] , 
       int_R_DATA_TEMPR123[8] ,int_R_DATA_TEMPR123[7] , 
       int_R_DATA_TEMPR123[6] ,int_R_DATA_TEMPR123[5] , 
       int_R_DATA_TEMPR123[4] ,int_R_DATA_TEMPR123[3] , 
       int_R_DATA_TEMPR123[2] ,int_R_DATA_TEMPR123[1] , 
       int_R_DATA_TEMPR123[0] }), .DB_DETECT(int_DB_DETECT_NG[123] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[123] ), .ACCESS_BUSY(
        ACCESS_BUSY[123] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[30] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[30] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR2 OR2_29 (.A(sel_R_DATA_TEMPR84[26] ), .B(sel_R_DATA_TEMPR85[26] ), .Y(
        OR2_29_Y));
    OR4 OR4_832 (.A(OR4_1303_Y), .B(OR4_1026_Y), .C(OR4_997_Y), .D(
        OR4_474_Y), .Y(OR4_832_Y));
    OR4 OR4_1385 (.A(sel_R_DATA_TEMPR72[7] ), .B(sel_R_DATA_TEMPR73[7] ), .C(sel_R_DATA_TEMPR74[7] ), .D(sel_R_DATA_TEMPR75[7] ), .Y(OR4_1385_Y));
    OR4 OR4_264 (.A(\DB_DETECT[48] ), .B(\DB_DETECT[49] ), .C(
        \DB_DETECT[50] ), .D(\DB_DETECT[51] ), .Y(OR4_264_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%22%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R22C0 (.A_DOUT({
        nc48, nc49, nc50, nc51, nc52,int_R_DATA_TEMPR22[31] , 
       int_R_DATA_TEMPR22[30] ,int_R_DATA_TEMPR22[29] , 
       int_R_DATA_TEMPR22[28] ,int_R_DATA_TEMPR22[27] , 
       int_R_DATA_TEMPR22[26] ,int_R_DATA_TEMPR22[25] , 
       int_R_DATA_TEMPR22[24] ,int_R_DATA_TEMPR22[23] , 
       int_R_DATA_TEMPR22[22] ,int_R_DATA_TEMPR22[21] , 
       int_R_DATA_TEMPR22[20] ,int_R_DATA_TEMPR22[19] , 
       int_R_DATA_TEMPR22[18] ,int_R_DATA_TEMPR22[17] }), .B_DOUT({nc53, 
        nc54, nc55,int_R_DATA_TEMPR22[16] ,int_R_DATA_TEMPR22[15] , 
       int_R_DATA_TEMPR22[14] ,int_R_DATA_TEMPR22[13] , 
       int_R_DATA_TEMPR22[12] ,int_R_DATA_TEMPR22[11] , 
       int_R_DATA_TEMPR22[10] ,int_R_DATA_TEMPR22[9] ,int_R_DATA_TEMPR22[8] , 
       int_R_DATA_TEMPR22[7] ,int_R_DATA_TEMPR22[6] ,int_R_DATA_TEMPR22[5] , 
       int_R_DATA_TEMPR22[4] ,int_R_DATA_TEMPR22[3] ,int_R_DATA_TEMPR22[2] , 
       int_R_DATA_TEMPR22[1] ,int_R_DATA_TEMPR22[0] }), .DB_DETECT( int_DB_DETECT_NG[22] ), .SB_CORRECT(int_SB_CORRECT_NG[22] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[22] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[5] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1340 (.A(sel_R_DATA_TEMPR88[24] ), .B(sel_R_DATA_TEMPR89[24] ), 
        .C(sel_R_DATA_TEMPR90[24] ), .D(sel_R_DATA_TEMPR91[24] ), .Y(
        OR4_1340_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%115%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R115C0 (.A_DOUT({
        nc56, nc57, nc58, nc59, nc60,int_R_DATA_TEMPR115[31] , 
       int_R_DATA_TEMPR115[30] ,int_R_DATA_TEMPR115[29] , 
       int_R_DATA_TEMPR115[28] ,int_R_DATA_TEMPR115[27] , 
       int_R_DATA_TEMPR115[26] ,int_R_DATA_TEMPR115[25] , 
       int_R_DATA_TEMPR115[24] ,int_R_DATA_TEMPR115[23] , 
       int_R_DATA_TEMPR115[22] ,int_R_DATA_TEMPR115[21] , 
       int_R_DATA_TEMPR115[20] ,int_R_DATA_TEMPR115[19] , 
       int_R_DATA_TEMPR115[18] ,int_R_DATA_TEMPR115[17] }), .B_DOUT({nc61, 
        nc62, nc63,int_R_DATA_TEMPR115[16] ,int_R_DATA_TEMPR115[15] , 
       int_R_DATA_TEMPR115[14] ,int_R_DATA_TEMPR115[13] , 
       int_R_DATA_TEMPR115[12] ,int_R_DATA_TEMPR115[11] , 
       int_R_DATA_TEMPR115[10] ,int_R_DATA_TEMPR115[9] , 
       int_R_DATA_TEMPR115[8] ,int_R_DATA_TEMPR115[7] , 
       int_R_DATA_TEMPR115[6] ,int_R_DATA_TEMPR115[5] , 
       int_R_DATA_TEMPR115[4] ,int_R_DATA_TEMPR115[3] , 
       int_R_DATA_TEMPR115[2] ,int_R_DATA_TEMPR115[1] , 
       int_R_DATA_TEMPR115[0] }), .DB_DETECT(int_DB_DETECT_NG[115] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[115] ), .ACCESS_BUSY(
        ACCESS_BUSY[115] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[28] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[28] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_656 (.A(\SB_CORRECT[88] ), .B(\SB_CORRECT[89] ), .C(
        \SB_CORRECT[90] ), .D(\SB_CORRECT[91] ), .Y(OR4_656_Y));
    OR4 OR4_1117 (.A(sel_R_DATA_TEMPR120[12] ), .B(sel_R_DATA_TEMPR121[12] ), 
        .C(sel_R_DATA_TEMPR122[12] ), .D(sel_R_DATA_TEMPR123[12] ), .Y(
        OR4_1117_Y));
    OR4 OR4_440 (.A(sel_R_DATA_TEMPR40[11] ), .B(sel_R_DATA_TEMPR41[11] ), 
        .C(sel_R_DATA_TEMPR42[11] ), .D(sel_R_DATA_TEMPR43[11] ), .Y(
        OR4_440_Y));
    AND4 \AND4DB_DETECT[22]  (.A(sel_DB_DETECT_NG[22] ), .B(
        \BLKY2_pipe[5] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[22] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%88%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R88C0 (.A_DOUT({
        nc64, nc65, nc66, nc67, nc68,int_R_DATA_TEMPR88[31] , 
       int_R_DATA_TEMPR88[30] ,int_R_DATA_TEMPR88[29] , 
       int_R_DATA_TEMPR88[28] ,int_R_DATA_TEMPR88[27] , 
       int_R_DATA_TEMPR88[26] ,int_R_DATA_TEMPR88[25] , 
       int_R_DATA_TEMPR88[24] ,int_R_DATA_TEMPR88[23] , 
       int_R_DATA_TEMPR88[22] ,int_R_DATA_TEMPR88[21] , 
       int_R_DATA_TEMPR88[20] ,int_R_DATA_TEMPR88[19] , 
       int_R_DATA_TEMPR88[18] ,int_R_DATA_TEMPR88[17] }), .B_DOUT({nc69, 
        nc70, nc71,int_R_DATA_TEMPR88[16] ,int_R_DATA_TEMPR88[15] , 
       int_R_DATA_TEMPR88[14] ,int_R_DATA_TEMPR88[13] , 
       int_R_DATA_TEMPR88[12] ,int_R_DATA_TEMPR88[11] , 
       int_R_DATA_TEMPR88[10] ,int_R_DATA_TEMPR88[9] ,int_R_DATA_TEMPR88[8] , 
       int_R_DATA_TEMPR88[7] ,int_R_DATA_TEMPR88[6] ,int_R_DATA_TEMPR88[5] , 
       int_R_DATA_TEMPR88[4] ,int_R_DATA_TEMPR88[3] ,int_R_DATA_TEMPR88[2] , 
       int_R_DATA_TEMPR88[1] ,int_R_DATA_TEMPR88[0] }), .DB_DETECT( int_DB_DETECT_NG[88] ), .SB_CORRECT(int_SB_CORRECT_NG[88] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[88] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[22] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4SB_CORRECT[0]  (.A(sel_SB_CORRECT_NG[0] ), .B(
        \BLKY2_pipe[0] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[0] ));
    OR4 OR4_1266 (.A(sel_R_DATA_TEMPR112[0] ), .B(sel_R_DATA_TEMPR113[0] ), 
        .C(sel_R_DATA_TEMPR114[0] ), .D(sel_R_DATA_TEMPR115[0] ), .Y(
        OR4_1266_Y));
    OR4 OR4_293 (.A(sel_R_DATA_TEMPR76[24] ), .B(sel_R_DATA_TEMPR77[24] ), 
        .C(sel_R_DATA_TEMPR78[24] ), .D(sel_R_DATA_TEMPR79[24] ), .Y(
        OR4_293_Y));
    OR4 OR4_388 (.A(OR4_980_Y), .B(OR4_835_Y), .C(OR4_947_Y), .D(
        OR4_974_Y), .Y(OR4_388_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%85%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R85C0 (.A_DOUT({
        nc72, nc73, nc74, nc75, nc76,int_R_DATA_TEMPR85[31] , 
       int_R_DATA_TEMPR85[30] ,int_R_DATA_TEMPR85[29] , 
       int_R_DATA_TEMPR85[28] ,int_R_DATA_TEMPR85[27] , 
       int_R_DATA_TEMPR85[26] ,int_R_DATA_TEMPR85[25] , 
       int_R_DATA_TEMPR85[24] ,int_R_DATA_TEMPR85[23] , 
       int_R_DATA_TEMPR85[22] ,int_R_DATA_TEMPR85[21] , 
       int_R_DATA_TEMPR85[20] ,int_R_DATA_TEMPR85[19] , 
       int_R_DATA_TEMPR85[18] ,int_R_DATA_TEMPR85[17] }), .B_DOUT({nc77, 
        nc78, nc79,int_R_DATA_TEMPR85[16] ,int_R_DATA_TEMPR85[15] , 
       int_R_DATA_TEMPR85[14] ,int_R_DATA_TEMPR85[13] , 
       int_R_DATA_TEMPR85[12] ,int_R_DATA_TEMPR85[11] , 
       int_R_DATA_TEMPR85[10] ,int_R_DATA_TEMPR85[9] ,int_R_DATA_TEMPR85[8] , 
       int_R_DATA_TEMPR85[7] ,int_R_DATA_TEMPR85[6] ,int_R_DATA_TEMPR85[5] , 
       int_R_DATA_TEMPR85[4] ,int_R_DATA_TEMPR85[3] ,int_R_DATA_TEMPR85[2] , 
       int_R_DATA_TEMPR85[1] ,int_R_DATA_TEMPR85[0] }), .DB_DETECT( int_DB_DETECT_NG[85] ), .SB_CORRECT(int_SB_CORRECT_NG[85] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[85] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[21] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[21] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_115 (.A(sel_R_DATA_TEMPR68[14] ), .B(sel_R_DATA_TEMPR69[14] ), 
        .C(sel_R_DATA_TEMPR70[14] ), .D(sel_R_DATA_TEMPR71[14] ), .Y(
        OR4_115_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%9%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R9C0 (.A_DOUT({
        nc80, nc81, nc82, nc83, nc84,int_R_DATA_TEMPR9[31] , 
       int_R_DATA_TEMPR9[30] ,int_R_DATA_TEMPR9[29] ,int_R_DATA_TEMPR9[28] , 
       int_R_DATA_TEMPR9[27] ,int_R_DATA_TEMPR9[26] ,int_R_DATA_TEMPR9[25] , 
       int_R_DATA_TEMPR9[24] ,int_R_DATA_TEMPR9[23] ,int_R_DATA_TEMPR9[22] , 
       int_R_DATA_TEMPR9[21] ,int_R_DATA_TEMPR9[20] ,int_R_DATA_TEMPR9[19] , 
       int_R_DATA_TEMPR9[18] ,int_R_DATA_TEMPR9[17] }), .B_DOUT({nc85, 
        nc86, nc87,int_R_DATA_TEMPR9[16] ,int_R_DATA_TEMPR9[15] , 
       int_R_DATA_TEMPR9[14] ,int_R_DATA_TEMPR9[13] ,int_R_DATA_TEMPR9[12] , 
       int_R_DATA_TEMPR9[11] ,int_R_DATA_TEMPR9[10] ,int_R_DATA_TEMPR9[9] , 
       int_R_DATA_TEMPR9[8] ,int_R_DATA_TEMPR9[7] ,int_R_DATA_TEMPR9[6] , 
       int_R_DATA_TEMPR9[5] ,int_R_DATA_TEMPR9[4] ,int_R_DATA_TEMPR9[3] , 
       int_R_DATA_TEMPR9[2] ,int_R_DATA_TEMPR9[1] ,int_R_DATA_TEMPR9[0] }), 
        .DB_DETECT(int_DB_DETECT_NG[9] ), .SB_CORRECT( int_SB_CORRECT_NG[9] ), .ACCESS_BUSY(\ACCESS_BUSY[9] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[2] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[2] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_66 (.A(sel_R_DATA_TEMPR52[7] ), .B(sel_R_DATA_TEMPR53[7] ), .C(sel_R_DATA_TEMPR54[7] ), .D(sel_R_DATA_TEMPR55[7] ), .Y(OR4_66_Y));
    OR4 OR4_1368 (.A(sel_R_DATA_TEMPR16[7] ), .B(sel_R_DATA_TEMPR17[7] ), .C(sel_R_DATA_TEMPR18[7] ), .D(sel_R_DATA_TEMPR19[7] ), .Y(OR4_1368_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[24]  (.A(CFG3_13_Y), .B(
        CFG3_7_Y), .Y(\BLKX2[24] ));
    OR4 OR4_998 (.A(sel_R_DATA_TEMPR28[31] ), .B(sel_R_DATA_TEMPR29[31] ), 
        .C(sel_R_DATA_TEMPR30[31] ), .D(sel_R_DATA_TEMPR31[31] ), .Y(
        OR4_998_Y));
    OR4 OR4_433 (.A(sel_R_DATA_TEMPR36[17] ), .B(sel_R_DATA_TEMPR37[17] ), 
        .C(sel_R_DATA_TEMPR38[17] ), .D(sel_R_DATA_TEMPR39[17] ), .Y(
        OR4_433_Y));
    OR4 OR4_417 (.A(OR4_1207_Y), .B(OR4_197_Y), .C(OR4_1012_Y), .D(
        OR4_1283_Y), .Y(OR4_417_Y));
    OR4 OR4_631 (.A(sel_R_DATA_TEMPR124[19] ), .B(sel_R_DATA_TEMPR125[19] ), 
        .C(sel_R_DATA_TEMPR126[19] ), .D(sel_R_DATA_TEMPR127[19] ), .Y(
        OR4_631_Y));
    OR4 OR4_365 (.A(sel_R_DATA_TEMPR44[5] ), .B(sel_R_DATA_TEMPR45[5] ), .C(sel_R_DATA_TEMPR46[5] ), .D(sel_R_DATA_TEMPR47[5] ), .Y(OR4_365_Y));
    OR4 OR4_238 (.A(sel_R_DATA_TEMPR100[4] ), .B(sel_R_DATA_TEMPR101[4] ), 
        .C(sel_R_DATA_TEMPR102[4] ), .D(sel_R_DATA_TEMPR103[4] ), .Y(
        OR4_238_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%61%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R61C0 (.A_DOUT({
        nc88, nc89, nc90, nc91, nc92,int_R_DATA_TEMPR61[31] , 
       int_R_DATA_TEMPR61[30] ,int_R_DATA_TEMPR61[29] , 
       int_R_DATA_TEMPR61[28] ,int_R_DATA_TEMPR61[27] , 
       int_R_DATA_TEMPR61[26] ,int_R_DATA_TEMPR61[25] , 
       int_R_DATA_TEMPR61[24] ,int_R_DATA_TEMPR61[23] , 
       int_R_DATA_TEMPR61[22] ,int_R_DATA_TEMPR61[21] , 
       int_R_DATA_TEMPR61[20] ,int_R_DATA_TEMPR61[19] , 
       int_R_DATA_TEMPR61[18] ,int_R_DATA_TEMPR61[17] }), .B_DOUT({nc93, 
        nc94, nc95,int_R_DATA_TEMPR61[16] ,int_R_DATA_TEMPR61[15] , 
       int_R_DATA_TEMPR61[14] ,int_R_DATA_TEMPR61[13] , 
       int_R_DATA_TEMPR61[12] ,int_R_DATA_TEMPR61[11] , 
       int_R_DATA_TEMPR61[10] ,int_R_DATA_TEMPR61[9] ,int_R_DATA_TEMPR61[8] , 
       int_R_DATA_TEMPR61[7] ,int_R_DATA_TEMPR61[6] ,int_R_DATA_TEMPR61[5] , 
       int_R_DATA_TEMPR61[4] ,int_R_DATA_TEMPR61[3] ,int_R_DATA_TEMPR61[2] , 
       int_R_DATA_TEMPR61[1] ,int_R_DATA_TEMPR61[0] }), .DB_DETECT( int_DB_DETECT_NG[61] ), .SB_CORRECT(int_SB_CORRECT_NG[61] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[61] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[15] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%90%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R90C0 (.A_DOUT({
        nc96, nc97, nc98, nc99, nc100,int_R_DATA_TEMPR90[31] , 
       int_R_DATA_TEMPR90[30] ,int_R_DATA_TEMPR90[29] , 
       int_R_DATA_TEMPR90[28] ,int_R_DATA_TEMPR90[27] , 
       int_R_DATA_TEMPR90[26] ,int_R_DATA_TEMPR90[25] , 
       int_R_DATA_TEMPR90[24] ,int_R_DATA_TEMPR90[23] , 
       int_R_DATA_TEMPR90[22] ,int_R_DATA_TEMPR90[21] , 
       int_R_DATA_TEMPR90[20] ,int_R_DATA_TEMPR90[19] , 
       int_R_DATA_TEMPR90[18] ,int_R_DATA_TEMPR90[17] }), .B_DOUT({nc101, 
        nc102, nc103,int_R_DATA_TEMPR90[16] ,int_R_DATA_TEMPR90[15] , 
       int_R_DATA_TEMPR90[14] ,int_R_DATA_TEMPR90[13] , 
       int_R_DATA_TEMPR90[12] ,int_R_DATA_TEMPR90[11] , 
       int_R_DATA_TEMPR90[10] ,int_R_DATA_TEMPR90[9] ,int_R_DATA_TEMPR90[8] , 
       int_R_DATA_TEMPR90[7] ,int_R_DATA_TEMPR90[6] ,int_R_DATA_TEMPR90[5] , 
       int_R_DATA_TEMPR90[4] ,int_R_DATA_TEMPR90[3] ,int_R_DATA_TEMPR90[2] , 
       int_R_DATA_TEMPR90[1] ,int_R_DATA_TEMPR90[0] }), .DB_DETECT( int_DB_DETECT_NG[90] ), .SB_CORRECT(int_SB_CORRECT_NG[90] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[90] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[22] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[22] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR2 OR2_8 (.A(sel_R_DATA_TEMPR84[24] ), .B(sel_R_DATA_TEMPR85[24] ), .Y(
        OR2_8_Y));
    AND4 \AND4DB_DETECT[76]  (.A(sel_DB_DETECT_NG[76] ), .B(
        \BLKY2_pipe[19] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[76] ));
    DFN1E1 \DFN1E1BLKY2_pipe[29]  (.D(\BLKY2[29] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[29] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%106%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R106C0 (.A_DOUT({
        nc104, nc105, nc106, nc107, nc108,int_R_DATA_TEMPR106[31] , 
       int_R_DATA_TEMPR106[30] ,int_R_DATA_TEMPR106[29] , 
       int_R_DATA_TEMPR106[28] ,int_R_DATA_TEMPR106[27] , 
       int_R_DATA_TEMPR106[26] ,int_R_DATA_TEMPR106[25] , 
       int_R_DATA_TEMPR106[24] ,int_R_DATA_TEMPR106[23] , 
       int_R_DATA_TEMPR106[22] ,int_R_DATA_TEMPR106[21] , 
       int_R_DATA_TEMPR106[20] ,int_R_DATA_TEMPR106[19] , 
       int_R_DATA_TEMPR106[18] ,int_R_DATA_TEMPR106[17] }), .B_DOUT({nc109, 
        nc110, nc111,int_R_DATA_TEMPR106[16] ,int_R_DATA_TEMPR106[15] , 
       int_R_DATA_TEMPR106[14] ,int_R_DATA_TEMPR106[13] , 
       int_R_DATA_TEMPR106[12] ,int_R_DATA_TEMPR106[11] , 
       int_R_DATA_TEMPR106[10] ,int_R_DATA_TEMPR106[9] , 
       int_R_DATA_TEMPR106[8] ,int_R_DATA_TEMPR106[7] , 
       int_R_DATA_TEMPR106[6] ,int_R_DATA_TEMPR106[5] , 
       int_R_DATA_TEMPR106[4] ,int_R_DATA_TEMPR106[3] , 
       int_R_DATA_TEMPR106[2] ,int_R_DATA_TEMPR106[1] , 
       int_R_DATA_TEMPR106[0] }), .DB_DETECT(int_DB_DETECT_NG[106] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[106] ), .ACCESS_BUSY(
        ACCESS_BUSY[106] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[26] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[26] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_189 (.A(OR4_93_Y), .B(OR4_473_Y), .C(OR4_1293_Y), .D(
        OR4_165_Y), .Y(OR4_189_Y));
    AND4 \AND4DB_DETECT[71]  (.A(sel_DB_DETECT_NG[71] ), .B(
        \BLKY2_pipe[17] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[71] ));
    OR4 OR4_0 (.A(sel_R_DATA_TEMPR80[11] ), .B(sel_R_DATA_TEMPR81[11] ), .C(sel_R_DATA_TEMPR82[11] ), .D(sel_R_DATA_TEMPR83[11] ), .Y(OR4_0_Y));
    OR4 OR4_207 (.A(OR4_348_Y), .B(OR2_29_Y), .C(sel_R_DATA_TEMPR86[26] ), 
        .D(sel_R_DATA_TEMPR87[26] ), .Y(OR4_207_Y));
    OR4 OR4_215 (.A(sel_R_DATA_TEMPR48[28] ), .B(sel_R_DATA_TEMPR49[28] ), 
        .C(sel_R_DATA_TEMPR50[28] ), .D(sel_R_DATA_TEMPR51[28] ), .Y(
        OR4_215_Y));
    AND4 \AND4SB_CORRECT[109]  (.A(sel_SB_CORRECT_NG[109] ), .B(
        \BLKY2_pipe[27] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[109] ));
    OR4 OR4_1245 (.A(OR4_106_Y), .B(OR4_1071_Y), .C(OR4_1121_Y), .D(
        OR4_601_Y), .Y(OR4_1245_Y));
    OR4 OR4_107 (.A(sel_R_DATA_TEMPR120[11] ), .B(sel_R_DATA_TEMPR121[11] ), 
        .C(sel_R_DATA_TEMPR122[11] ), .D(sel_R_DATA_TEMPR123[11] ), .Y(
        OR4_107_Y));
    OR4 OR4_1002 (.A(\SB_CORRECT[48] ), .B(\SB_CORRECT[49] ), .C(
        \SB_CORRECT[50] ), .D(\SB_CORRECT[51] ), .Y(OR4_1002_Y));
    OR4 OR4_1069 (.A(sel_R_DATA_TEMPR4[11] ), .B(sel_R_DATA_TEMPR5[11] ), .C(sel_R_DATA_TEMPR6[11] ), .D(sel_R_DATA_TEMPR7[11] ), .Y(OR4_1069_Y));
    AND4 \AND4SB_CORRECT[28]  (.A(sel_SB_CORRECT_NG[28] ), .B(
        \BLKY2_pipe[7] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[28] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%39%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R39C0 (.A_DOUT({
        nc112, nc113, nc114, nc115, nc116,int_R_DATA_TEMPR39[31] , 
       int_R_DATA_TEMPR39[30] ,int_R_DATA_TEMPR39[29] , 
       int_R_DATA_TEMPR39[28] ,int_R_DATA_TEMPR39[27] , 
       int_R_DATA_TEMPR39[26] ,int_R_DATA_TEMPR39[25] , 
       int_R_DATA_TEMPR39[24] ,int_R_DATA_TEMPR39[23] , 
       int_R_DATA_TEMPR39[22] ,int_R_DATA_TEMPR39[21] , 
       int_R_DATA_TEMPR39[20] ,int_R_DATA_TEMPR39[19] , 
       int_R_DATA_TEMPR39[18] ,int_R_DATA_TEMPR39[17] }), .B_DOUT({nc117, 
        nc118, nc119,int_R_DATA_TEMPR39[16] ,int_R_DATA_TEMPR39[15] , 
       int_R_DATA_TEMPR39[14] ,int_R_DATA_TEMPR39[13] , 
       int_R_DATA_TEMPR39[12] ,int_R_DATA_TEMPR39[11] , 
       int_R_DATA_TEMPR39[10] ,int_R_DATA_TEMPR39[9] ,int_R_DATA_TEMPR39[8] , 
       int_R_DATA_TEMPR39[7] ,int_R_DATA_TEMPR39[6] ,int_R_DATA_TEMPR39[5] , 
       int_R_DATA_TEMPR39[4] ,int_R_DATA_TEMPR39[3] ,int_R_DATA_TEMPR39[2] , 
       int_R_DATA_TEMPR39[1] ,int_R_DATA_TEMPR39[0] }), .DB_DETECT( int_DB_DETECT_NG[39] ), .SB_CORRECT(int_SB_CORRECT_NG[39] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[39] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[9] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[9] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_812 (.A(sel_R_DATA_TEMPR92[24] ), .B(sel_R_DATA_TEMPR93[24] ), 
        .C(sel_R_DATA_TEMPR94[24] ), .D(sel_R_DATA_TEMPR95[24] ), .Y(
        OR4_812_Y));
    OR4 OR4_277 (.A(OR4_119_Y), .B(OR4_1298_Y), .C(OR4_1049_Y), .D(
        OR4_40_Y), .Y(OR4_277_Y));
    OR4 OR4_698 (.A(sel_R_DATA_TEMPR68[26] ), .B(sel_R_DATA_TEMPR69[26] ), 
        .C(sel_R_DATA_TEMPR70[26] ), .D(sel_R_DATA_TEMPR71[26] ), .Y(
        OR4_698_Y));
    OR4 OR4_95 (.A(sel_R_DATA_TEMPR44[3] ), .B(sel_R_DATA_TEMPR45[3] ), .C(sel_R_DATA_TEMPR46[3] ), .D(sel_R_DATA_TEMPR47[3] ), .Y(OR4_95_Y));
    OR2 OR2_22 (.A(\SB_CORRECT[84] ), .B(\SB_CORRECT[85] ), .Y(
        OR2_22_Y));
    OR4 OR4_177 (.A(sel_R_DATA_TEMPR80[20] ), .B(sel_R_DATA_TEMPR81[20] ), 
        .C(sel_R_DATA_TEMPR82[20] ), .D(sel_R_DATA_TEMPR83[20] ), .Y(
        OR4_177_Y));
    OR4 OR4_981 (.A(sel_R_DATA_TEMPR8[2] ), .B(sel_R_DATA_TEMPR9[2] ), .C(sel_R_DATA_TEMPR10[2] ), .D(sel_R_DATA_TEMPR11[2] ), .Y(OR4_981_Y));
    OR4 OR4_1296 (.A(sel_R_DATA_TEMPR124[7] ), .B(sel_R_DATA_TEMPR125[7] ), 
        .C(sel_R_DATA_TEMPR126[7] ), .D(sel_R_DATA_TEMPR127[7] ), .Y(
        OR4_1296_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[14]  (.A(CFG3_1_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[14] ));
    AND4 \AND4DB_DETECT[87]  (.A(sel_DB_DETECT_NG[87] ), .B(
        \BLKY2_pipe[21] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[87] ));
    OR4 OR4_762 (.A(OR4_808_Y), .B(OR2_10_Y), .C(\DB_DETECT[86] ), 
        .D(\DB_DETECT[87] ), .Y(OR4_762_Y));
    OR4 OR4_349 (.A(sel_R_DATA_TEMPR108[26] ), .B(sel_R_DATA_TEMPR109[26] ), 
        .C(sel_R_DATA_TEMPR110[26] ), .D(sel_R_DATA_TEMPR111[26] ), .Y(
        OR4_349_Y));
    OR4 OR4_1239 (.A(sel_R_DATA_TEMPR88[25] ), .B(sel_R_DATA_TEMPR89[25] ), 
        .C(sel_R_DATA_TEMPR90[25] ), .D(sel_R_DATA_TEMPR91[25] ), .Y(
        OR4_1239_Y));
    OR4 OR4_692 (.A(\DB_DETECT[116] ), .B(\DB_DETECT[117] ), .C(
        \DB_DETECT[118] ), .D(\DB_DETECT[119] ), .Y(OR4_692_Y));
    OR4 OR4_1210 (.A(sel_R_DATA_TEMPR4[10] ), .B(sel_R_DATA_TEMPR5[10] ), .C(sel_R_DATA_TEMPR6[10] ), .D(sel_R_DATA_TEMPR7[10] ), .Y(OR4_1210_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[31]  (.A(CFG3_21_Y), .B(
        CFG3_3_Y), .Y(\BLKY2[31] ));
    OR4 OR4_703 (.A(sel_R_DATA_TEMPR80[28] ), .B(sel_R_DATA_TEMPR81[28] ), 
        .C(sel_R_DATA_TEMPR82[28] ), .D(sel_R_DATA_TEMPR83[28] ), .Y(
        OR4_703_Y));
    OR4 OR4_223 (.A(OR4_621_Y), .B(OR4_1094_Y), .C(OR4_978_Y), .D(
        OR4_421_Y), .Y(OR4_223_Y));
    OR4 OR4_966 (.A(OR4_841_Y), .B(OR4_337_Y), .C(OR4_542_Y), .D(
        OR4_1034_Y), .Y(OR4_966_Y));
    OR4 OR4_204 (.A(sel_R_DATA_TEMPR60[28] ), .B(sel_R_DATA_TEMPR61[28] ), 
        .C(sel_R_DATA_TEMPR62[28] ), .D(sel_R_DATA_TEMPR63[28] ), .Y(
        OR4_204_Y));
    OR4 OR4_354 (.A(sel_R_DATA_TEMPR44[0] ), .B(sel_R_DATA_TEMPR45[0] ), .C(sel_R_DATA_TEMPR46[0] ), .D(sel_R_DATA_TEMPR47[0] ), .Y(OR4_354_Y));
    OR2 OR2_19 (.A(sel_R_DATA_TEMPR84[5] ), .B(sel_R_DATA_TEMPR85[5] ), .Y(
        OR2_19_Y));
    OR4 OR4_773 (.A(OR4_868_Y), .B(OR4_1102_Y), .C(OR4_673_Y), .D(
        OR4_466_Y), .Y(OR4_773_Y));
    OR4 OR4_665 (.A(sel_R_DATA_TEMPR8[27] ), .B(sel_R_DATA_TEMPR9[27] ), .C(sel_R_DATA_TEMPR10[27] ), .D(sel_R_DATA_TEMPR11[27] ), .Y(OR4_665_Y));
    OR4 OR4_413 (.A(sel_R_DATA_TEMPR88[18] ), .B(sel_R_DATA_TEMPR89[18] ), 
        .C(sel_R_DATA_TEMPR90[18] ), .D(sel_R_DATA_TEMPR91[18] ), .Y(
        OR4_413_Y));
    OR4 OR4_611 (.A(sel_R_DATA_TEMPR80[12] ), .B(sel_R_DATA_TEMPR81[12] ), 
        .C(sel_R_DATA_TEMPR82[12] ), .D(sel_R_DATA_TEMPR83[12] ), .Y(
        OR4_611_Y));
    OR4 OR4_1312 (.A(sel_R_DATA_TEMPR44[4] ), .B(sel_R_DATA_TEMPR45[4] ), .C(sel_R_DATA_TEMPR46[4] ), .D(sel_R_DATA_TEMPR47[4] ), .Y(OR4_1312_Y));
    OR4 OR4_1082 (.A(OR4_782_Y), .B(OR4_564_Y), .C(OR4_332_Y), .D(
        OR4_293_Y), .Y(OR4_1082_Y));
    OR4 OR4_928 (.A(sel_R_DATA_TEMPR28[23] ), .B(sel_R_DATA_TEMPR29[23] ), 
        .C(sel_R_DATA_TEMPR30[23] ), .D(sel_R_DATA_TEMPR31[23] ), .Y(
        OR4_928_Y));
    OR4 OR4_151 (.A(sel_R_DATA_TEMPR24[16] ), .B(sel_R_DATA_TEMPR25[16] ), 
        .C(sel_R_DATA_TEMPR26[16] ), .D(sel_R_DATA_TEMPR27[16] ), .Y(
        OR4_151_Y));
    OR4 OR4_274 (.A(OR4_823_Y), .B(OR4_685_Y), .C(OR4_786_Y), .D(
        OR4_651_Y), .Y(OR4_274_Y));
    AND4 \AND4DB_DETECT[39]  (.A(sel_DB_DETECT_NG[39] ), .B(
        \BLKY2_pipe[9] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[39] ));
    OR4 OR4_218 (.A(OR4_169_Y), .B(OR2_17_Y), .C(sel_R_DATA_TEMPR86[9] ), 
        .D(sel_R_DATA_TEMPR87[9] ), .Y(OR4_218_Y));
    OR4 OR4_1212 (.A(OR4_271_Y), .B(OR4_115_Y), .C(OR4_232_Y), .D(
        OR4_1242_Y), .Y(OR4_1212_Y));
    OR4 \OR4_R_DATA[22]  (.A(OR4_873_Y), .B(OR4_834_Y), .C(OR4_646_Y), 
        .D(OR4_31_Y), .Y(R_DATA[22]));
    OR4 OR4_60 (.A(sel_R_DATA_TEMPR40[29] ), .B(sel_R_DATA_TEMPR41[29] ), .C(sel_R_DATA_TEMPR42[29] ), .D(sel_R_DATA_TEMPR43[29] ), .Y(OR4_60_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%0%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R0C0 (.A_DOUT({
        nc120, nc121, nc122, nc123, nc124,int_R_DATA_TEMPR0[31] , 
       int_R_DATA_TEMPR0[30] ,int_R_DATA_TEMPR0[29] ,int_R_DATA_TEMPR0[28] , 
       int_R_DATA_TEMPR0[27] ,int_R_DATA_TEMPR0[26] ,int_R_DATA_TEMPR0[25] , 
       int_R_DATA_TEMPR0[24] ,int_R_DATA_TEMPR0[23] ,int_R_DATA_TEMPR0[22] , 
       int_R_DATA_TEMPR0[21] ,int_R_DATA_TEMPR0[20] ,int_R_DATA_TEMPR0[19] , 
       int_R_DATA_TEMPR0[18] ,int_R_DATA_TEMPR0[17] }), .B_DOUT({nc125, 
        nc126, nc127,int_R_DATA_TEMPR0[16] ,int_R_DATA_TEMPR0[15] , 
       int_R_DATA_TEMPR0[14] ,int_R_DATA_TEMPR0[13] ,int_R_DATA_TEMPR0[12] , 
       int_R_DATA_TEMPR0[11] ,int_R_DATA_TEMPR0[10] ,int_R_DATA_TEMPR0[9] , 
       int_R_DATA_TEMPR0[8] ,int_R_DATA_TEMPR0[7] ,int_R_DATA_TEMPR0[6] , 
       int_R_DATA_TEMPR0[5] ,int_R_DATA_TEMPR0[4] ,int_R_DATA_TEMPR0[3] , 
       int_R_DATA_TEMPR0[2] ,int_R_DATA_TEMPR0[1] ,int_R_DATA_TEMPR0[0] }), 
        .DB_DETECT(int_DB_DETECT_NG[0] ), .SB_CORRECT( int_SB_CORRECT_NG[0] ), .ACCESS_BUSY(\ACCESS_BUSY[0] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4SB_CORRECT[68]  (.A(sel_SB_CORRECT_NG[68] ), .B(
        \BLKY2_pipe[17] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[68] ));
    OR4 OR4_1355 (.A(OR4_849_Y), .B(OR2_3_Y), .C(sel_R_DATA_TEMPR86[13] ), 
        .D(sel_R_DATA_TEMPR87[13] ), .Y(OR4_1355_Y));
    AND4 \AND4SB_CORRECT[87]  (.A(sel_SB_CORRECT_NG[87] ), .B(
        \BLKY2_pipe[21] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[87] ));
    OR4 OR4_531 (.A(sel_R_DATA_TEMPR20[24] ), .B(sel_R_DATA_TEMPR21[24] ), 
        .C(sel_R_DATA_TEMPR22[24] ), .D(sel_R_DATA_TEMPR23[24] ), .Y(
        OR4_531_Y));
    OR4 OR4_1099 (.A(sel_R_DATA_TEMPR76[9] ), .B(sel_R_DATA_TEMPR77[9] ), .C(sel_R_DATA_TEMPR78[9] ), .D(sel_R_DATA_TEMPR79[9] ), .Y(OR4_1099_Y));
    OR4 OR4_895 (.A(sel_R_DATA_TEMPR36[21] ), .B(sel_R_DATA_TEMPR37[21] ), 
        .C(sel_R_DATA_TEMPR38[21] ), .D(sel_R_DATA_TEMPR39[21] ), .Y(
        OR4_895_Y));
    OR4 OR4_67 (.A(sel_R_DATA_TEMPR16[14] ), .B(sel_R_DATA_TEMPR17[14] ), .C(sel_R_DATA_TEMPR18[14] ), .D(sel_R_DATA_TEMPR19[14] ), .Y(OR4_67_Y));
    OR4 OR4_785 (.A(OR4_668_Y), .B(OR4_461_Y), .C(OR4_213_Y), .D(
        OR4_864_Y), .Y(OR4_785_Y));
    OR4 OR4_687 (.A(OR4_177_Y), .B(OR2_26_Y), .C(sel_R_DATA_TEMPR86[20] ), 
        .D(sel_R_DATA_TEMPR87[20] ), .Y(OR4_687_Y));
    OR4 OR4_305 (.A(OR4_1107_Y), .B(OR4_1373_Y), .C(OR4_889_Y), .D(
        OR4_237_Y), .Y(OR4_305_Y));
    OR4 OR4_451 (.A(sel_R_DATA_TEMPR12[7] ), .B(sel_R_DATA_TEMPR13[7] ), .C(sel_R_DATA_TEMPR14[7] ), .D(sel_R_DATA_TEMPR15[7] ), .Y(OR4_451_Y));
    OR4 OR4_1214 (.A(OR4_769_Y), .B(OR4_496_Y), .C(OR4_268_Y), .D(
        OR4_328_Y), .Y(OR4_1214_Y));
    OR4 OR4_786 (.A(sel_R_DATA_TEMPR72[10] ), .B(sel_R_DATA_TEMPR73[10] ), 
        .C(sel_R_DATA_TEMPR74[10] ), .D(sel_R_DATA_TEMPR75[10] ), .Y(
        OR4_786_Y));
    OR4 OR4_458 (.A(sel_R_DATA_TEMPR16[22] ), .B(sel_R_DATA_TEMPR17[22] ), 
        .C(sel_R_DATA_TEMPR18[22] ), .D(sel_R_DATA_TEMPR19[22] ), .Y(
        OR4_458_Y));
    OR4 OR4_1173 (.A(sel_R_DATA_TEMPR80[7] ), .B(sel_R_DATA_TEMPR81[7] ), .C(sel_R_DATA_TEMPR82[7] ), .D(sel_R_DATA_TEMPR83[7] ), .Y(OR4_1173_Y));
    OR4 OR4_628 (.A(sel_R_DATA_TEMPR96[3] ), .B(sel_R_DATA_TEMPR97[3] ), .C(sel_R_DATA_TEMPR98[3] ), .D(sel_R_DATA_TEMPR99[3] ), .Y(OR4_628_Y));
    OR4 OR4_375 (.A(sel_R_DATA_TEMPR68[30] ), .B(sel_R_DATA_TEMPR69[30] ), 
        .C(sel_R_DATA_TEMPR70[30] ), .D(sel_R_DATA_TEMPR71[30] ), .Y(
        OR4_375_Y));
    OR4 OR4_1317 (.A(\DB_DETECT[16] ), .B(\DB_DETECT[17] ), .C(
        \DB_DETECT[18] ), .D(\DB_DETECT[19] ), .Y(OR4_1317_Y));
    OR4 OR4_749 (.A(sel_R_DATA_TEMPR20[5] ), .B(sel_R_DATA_TEMPR21[5] ), .C(sel_R_DATA_TEMPR22[5] ), .D(sel_R_DATA_TEMPR23[5] ), .Y(OR4_749_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%47%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R47C0 (.A_DOUT({
        nc128, nc129, nc130, nc131, nc132,int_R_DATA_TEMPR47[31] , 
       int_R_DATA_TEMPR47[30] ,int_R_DATA_TEMPR47[29] , 
       int_R_DATA_TEMPR47[28] ,int_R_DATA_TEMPR47[27] , 
       int_R_DATA_TEMPR47[26] ,int_R_DATA_TEMPR47[25] , 
       int_R_DATA_TEMPR47[24] ,int_R_DATA_TEMPR47[23] , 
       int_R_DATA_TEMPR47[22] ,int_R_DATA_TEMPR47[21] , 
       int_R_DATA_TEMPR47[20] ,int_R_DATA_TEMPR47[19] , 
       int_R_DATA_TEMPR47[18] ,int_R_DATA_TEMPR47[17] }), .B_DOUT({nc133, 
        nc134, nc135,int_R_DATA_TEMPR47[16] ,int_R_DATA_TEMPR47[15] , 
       int_R_DATA_TEMPR47[14] ,int_R_DATA_TEMPR47[13] , 
       int_R_DATA_TEMPR47[12] ,int_R_DATA_TEMPR47[11] , 
       int_R_DATA_TEMPR47[10] ,int_R_DATA_TEMPR47[9] ,int_R_DATA_TEMPR47[8] , 
       int_R_DATA_TEMPR47[7] ,int_R_DATA_TEMPR47[6] ,int_R_DATA_TEMPR47[5] , 
       int_R_DATA_TEMPR47[4] ,int_R_DATA_TEMPR47[3] ,int_R_DATA_TEMPR47[2] , 
       int_R_DATA_TEMPR47[1] ,int_R_DATA_TEMPR47[0] }), .DB_DETECT( int_DB_DETECT_NG[47] ), .SB_CORRECT(int_SB_CORRECT_NG[47] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[47] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[11] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[11] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1229 (.A(OR4_532_Y), .B(OR4_1270_Y), .C(OR4_551_Y), .D(
        OR4_763_Y), .Y(OR4_1229_Y));
    OR4 OR4_660 (.A(OR4_247_Y), .B(OR4_538_Y), .C(OR4_515_Y), .D(
        OR4_1190_Y), .Y(OR4_660_Y));
    AND4 \AND4DB_DETECT[10]  (.A(sel_DB_DETECT_NG[10] ), .B(
        \BLKY2_pipe[2] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[10] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%23%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R23C0 (.A_DOUT({
        nc136, nc137, nc138, nc139, nc140,int_R_DATA_TEMPR23[31] , 
       int_R_DATA_TEMPR23[30] ,int_R_DATA_TEMPR23[29] , 
       int_R_DATA_TEMPR23[28] ,int_R_DATA_TEMPR23[27] , 
       int_R_DATA_TEMPR23[26] ,int_R_DATA_TEMPR23[25] , 
       int_R_DATA_TEMPR23[24] ,int_R_DATA_TEMPR23[23] , 
       int_R_DATA_TEMPR23[22] ,int_R_DATA_TEMPR23[21] , 
       int_R_DATA_TEMPR23[20] ,int_R_DATA_TEMPR23[19] , 
       int_R_DATA_TEMPR23[18] ,int_R_DATA_TEMPR23[17] }), .B_DOUT({nc141, 
        nc142, nc143,int_R_DATA_TEMPR23[16] ,int_R_DATA_TEMPR23[15] , 
       int_R_DATA_TEMPR23[14] ,int_R_DATA_TEMPR23[13] , 
       int_R_DATA_TEMPR23[12] ,int_R_DATA_TEMPR23[11] , 
       int_R_DATA_TEMPR23[10] ,int_R_DATA_TEMPR23[9] ,int_R_DATA_TEMPR23[8] , 
       int_R_DATA_TEMPR23[7] ,int_R_DATA_TEMPR23[6] ,int_R_DATA_TEMPR23[5] , 
       int_R_DATA_TEMPR23[4] ,int_R_DATA_TEMPR23[3] ,int_R_DATA_TEMPR23[2] , 
       int_R_DATA_TEMPR23[1] ,int_R_DATA_TEMPR23[0] }), .DB_DETECT( int_DB_DETECT_NG[23] ), .SB_CORRECT(int_SB_CORRECT_NG[23] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[23] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[5] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_622 (.A(sel_R_DATA_TEMPR16[16] ), .B(sel_R_DATA_TEMPR17[16] ), 
        .C(sel_R_DATA_TEMPR18[16] ), .D(sel_R_DATA_TEMPR19[16] ), .Y(
        OR4_622_Y));
    OR4 OR4_232 (.A(sel_R_DATA_TEMPR72[14] ), .B(sel_R_DATA_TEMPR73[14] ), 
        .C(sel_R_DATA_TEMPR74[14] ), .D(sel_R_DATA_TEMPR75[14] ), .Y(
        OR4_232_Y));
    OR4 OR4_844 (.A(sel_R_DATA_TEMPR120[26] ), .B(sel_R_DATA_TEMPR121[26] ), 
        .C(sel_R_DATA_TEMPR122[26] ), .D(sel_R_DATA_TEMPR123[26] ), .Y(
        OR4_844_Y));
    AND4 \AND4SB_CORRECT[5]  (.A(sel_SB_CORRECT_NG[5] ), .B(
        \BLKY2_pipe[1] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[5] ));
    CFG3 #( .INIT(8'h2) )  CFG3_6 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_6_Y));
    OR4 \OR4_R_DATA[15]  (.A(OR4_1218_Y), .B(OR4_485_Y), .C(OR4_1011_Y)
        , .D(OR4_618_Y), .Y(R_DATA[15]));
    OR4 OR4_1167 (.A(sel_R_DATA_TEMPR76[0] ), .B(sel_R_DATA_TEMPR77[0] ), .C(sel_R_DATA_TEMPR78[0] ), .D(sel_R_DATA_TEMPR79[0] ), .Y(OR4_1167_Y));
    OR4 OR4_543 (.A(OR4_1169_Y), .B(OR4_45_Y), .C(OR4_251_Y), .D(
        OR4_92_Y), .Y(OR4_543_Y));
    OR2 OR2_12 (.A(sel_R_DATA_TEMPR84[18] ), .B(sel_R_DATA_TEMPR85[18] ), .Y(
        OR2_12_Y));
    DFN1E1 \DFN1E1BLKY1_pipe[0]  (.D(\BLKY1[0] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY1_pipe[0] ));
    OR4 OR4_45 (.A(sel_R_DATA_TEMPR52[15] ), .B(sel_R_DATA_TEMPR53[15] ), .C(sel_R_DATA_TEMPR54[15] ), .D(sel_R_DATA_TEMPR55[15] ), .Y(OR4_45_Y));
    OR4 OR4_367 (.A(OR4_1223_Y), .B(OR4_757_Y), .C(OR4_1239_Y), .D(
        OR4_704_Y), .Y(OR4_367_Y));
    OR4 OR4_160 (.A(OR4_746_Y), .B(OR4_1134_Y), .C(OR4_563_Y), .D(
        OR4_821_Y), .Y(OR4_160_Y));
    OR4 OR4_702 (.A(sel_R_DATA_TEMPR60[16] ), .B(sel_R_DATA_TEMPR61[16] ), 
        .C(sel_R_DATA_TEMPR62[16] ), .D(sel_R_DATA_TEMPR63[16] ), .Y(
        OR4_702_Y));
    OR4 OR4_559 (.A(OR4_164_Y), .B(OR2_25_Y), .C(sel_R_DATA_TEMPR86[22] ), 
        .D(sel_R_DATA_TEMPR87[22] ), .Y(OR4_559_Y));
    AND4 \AND4SB_CORRECT[41]  (.A(sel_SB_CORRECT_NG[41] ), .B(
        \BLKY2_pipe[10] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[41] ));
    OR4 OR4_1044 (.A(sel_R_DATA_TEMPR100[23] ), .B(sel_R_DATA_TEMPR101[23] ), 
        .C(sel_R_DATA_TEMPR102[23] ), .D(sel_R_DATA_TEMPR103[23] ), .Y(
        OR4_1044_Y));
    OR4 OR4_550 (.A(sel_R_DATA_TEMPR76[17] ), .B(sel_R_DATA_TEMPR77[17] ), 
        .C(sel_R_DATA_TEMPR78[17] ), .D(sel_R_DATA_TEMPR79[17] ), .Y(
        OR4_550_Y));
    OR4 \OR4_R_DATA[23]  (.A(OR4_723_Y), .B(OR4_368_Y), .C(OR4_313_Y), 
        .D(OR4_277_Y), .Y(R_DATA[23]));
    OR4 OR4_330 (.A(OR4_352_Y), .B(OR4_604_Y), .C(OR4_138_Y), .D(
        OR4_855_Y), .Y(OR4_330_Y));
    OR4 OR4_906 (.A(OR4_1189_Y), .B(OR4_976_Y), .C(OR4_58_Y), .D(
        OR4_446_Y), .Y(OR4_906_Y));
    OR4 OR4_772 (.A(OR4_143_Y), .B(OR2_15_Y), .C(sel_R_DATA_TEMPR86[2] ), 
        .D(sel_R_DATA_TEMPR87[2] ), .Y(OR4_772_Y));
    OR4 OR4_768 (.A(sel_R_DATA_TEMPR4[1] ), .B(sel_R_DATA_TEMPR5[1] ), .C(sel_R_DATA_TEMPR6[1] ), .D(sel_R_DATA_TEMPR7[1] ), .Y(OR4_768_Y));
    OR4 OR4_1343 (.A(sel_R_DATA_TEMPR88[28] ), .B(sel_R_DATA_TEMPR89[28] ), 
        .C(sel_R_DATA_TEMPR90[28] ), .D(sel_R_DATA_TEMPR91[28] ), .Y(
        OR4_1343_Y));
    AND4 \AND4SB_CORRECT[118]  (.A(sel_SB_CORRECT_NG[118] ), .B(
        \BLKY2_pipe[29] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[118] ));
    OR4 OR4_605 (.A(sel_R_DATA_TEMPR0[19] ), .B(sel_R_DATA_TEMPR1[19] ), .C(sel_R_DATA_TEMPR2[19] ), .D(sel_R_DATA_TEMPR3[19] ), .Y(OR4_605_Y));
    OR4 OR4_511 (.A(sel_R_DATA_TEMPR28[20] ), .B(sel_R_DATA_TEMPR29[20] ), 
        .C(sel_R_DATA_TEMPR30[20] ), .D(sel_R_DATA_TEMPR31[20] ), .Y(
        OR4_511_Y));
    OR4 OR4_976 (.A(sel_R_DATA_TEMPR36[2] ), .B(sel_R_DATA_TEMPR37[2] ), .C(sel_R_DATA_TEMPR38[2] ), .D(sel_R_DATA_TEMPR39[2] ), .Y(OR4_976_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[20]  (.A(CFG3_6_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[20] ));
    OR4 OR4_1233 (.A(sel_R_DATA_TEMPR60[12] ), .B(sel_R_DATA_TEMPR61[12] ), 
        .C(sel_R_DATA_TEMPR62[12] ), .D(sel_R_DATA_TEMPR63[12] ), .Y(
        OR4_1233_Y));
    OR4 OR4_833 (.A(sel_R_DATA_TEMPR68[8] ), .B(sel_R_DATA_TEMPR69[8] ), .C(sel_R_DATA_TEMPR70[8] ), .D(sel_R_DATA_TEMPR71[8] ), .Y(OR4_833_Y));
    OR4 OR4_825 (.A(sel_R_DATA_TEMPR28[14] ), .B(sel_R_DATA_TEMPR29[14] ), 
        .C(sel_R_DATA_TEMPR30[14] ), .D(sel_R_DATA_TEMPR31[14] ), .Y(
        OR4_825_Y));
    OR4 OR4_696 (.A(sel_R_DATA_TEMPR108[22] ), .B(sel_R_DATA_TEMPR109[22] ), 
        .C(sel_R_DATA_TEMPR110[22] ), .D(sel_R_DATA_TEMPR111[22] ), .Y(
        OR4_696_Y));
    OR4 OR4_675 (.A(sel_R_DATA_TEMPR12[25] ), .B(sel_R_DATA_TEMPR13[25] ), 
        .C(sel_R_DATA_TEMPR14[25] ), .D(sel_R_DATA_TEMPR15[25] ), .Y(
        OR4_675_Y));
    OR4 OR4_287 (.A(sel_R_DATA_TEMPR80[19] ), .B(sel_R_DATA_TEMPR81[19] ), 
        .C(sel_R_DATA_TEMPR82[19] ), .D(sel_R_DATA_TEMPR83[19] ), .Y(
        OR4_287_Y));
    OR4 OR4_86 (.A(sel_R_DATA_TEMPR36[6] ), .B(sel_R_DATA_TEMPR37[6] ), .C(sel_R_DATA_TEMPR38[6] ), .D(sel_R_DATA_TEMPR39[6] ), .Y(OR4_86_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%5%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R5C0 (.A_DOUT({
        nc144, nc145, nc146, nc147, nc148,int_R_DATA_TEMPR5[31] , 
       int_R_DATA_TEMPR5[30] ,int_R_DATA_TEMPR5[29] ,int_R_DATA_TEMPR5[28] , 
       int_R_DATA_TEMPR5[27] ,int_R_DATA_TEMPR5[26] ,int_R_DATA_TEMPR5[25] , 
       int_R_DATA_TEMPR5[24] ,int_R_DATA_TEMPR5[23] ,int_R_DATA_TEMPR5[22] , 
       int_R_DATA_TEMPR5[21] ,int_R_DATA_TEMPR5[20] ,int_R_DATA_TEMPR5[19] , 
       int_R_DATA_TEMPR5[18] ,int_R_DATA_TEMPR5[17] }), .B_DOUT({nc149, 
        nc150, nc151,int_R_DATA_TEMPR5[16] ,int_R_DATA_TEMPR5[15] , 
       int_R_DATA_TEMPR5[14] ,int_R_DATA_TEMPR5[13] ,int_R_DATA_TEMPR5[12] , 
       int_R_DATA_TEMPR5[11] ,int_R_DATA_TEMPR5[10] ,int_R_DATA_TEMPR5[9] , 
       int_R_DATA_TEMPR5[8] ,int_R_DATA_TEMPR5[7] ,int_R_DATA_TEMPR5[6] , 
       int_R_DATA_TEMPR5[5] ,int_R_DATA_TEMPR5[4] ,int_R_DATA_TEMPR5[3] , 
       int_R_DATA_TEMPR5[2] ,int_R_DATA_TEMPR5[1] ,int_R_DATA_TEMPR5[0] }), 
        .DB_DETECT(int_DB_DETECT_NG[5] ), .SB_CORRECT( int_SB_CORRECT_NG[5] ), .ACCESS_BUSY(\ACCESS_BUSY[5] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[4]  (.A(CFG3_6_Y), .B(CFG3_12_Y)
        , .Y(\BLKX2[4] ));
    OR4 OR4_33 (.A(sel_R_DATA_TEMPR12[8] ), .B(sel_R_DATA_TEMPR13[8] ), .C(sel_R_DATA_TEMPR14[8] ), .D(sel_R_DATA_TEMPR15[8] ), .Y(OR4_33_Y));
    AND4 \AND4DB_DETECT[108]  (.A(sel_DB_DETECT_NG[108] ), .B(
        \BLKY2_pipe[27] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[108] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[10]  (.A(CFG3_0_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[10] ));
    OR4 OR4_867 (.A(OR4_152_Y), .B(OR4_1027_Y), .C(OR4_1248_Y), .D(
        OR4_340_Y), .Y(OR4_867_Y));
    OR4 OR4_168 (.A(OR4_754_Y), .B(OR4_480_Y), .C(OR4_923_Y), .D(
        OR4_1312_Y), .Y(OR4_168_Y));
    OR4 OR4_964 (.A(sel_R_DATA_TEMPR24[14] ), .B(sel_R_DATA_TEMPR25[14] ), 
        .C(sel_R_DATA_TEMPR26[14] ), .D(sel_R_DATA_TEMPR27[14] ), .Y(
        OR4_964_Y));
    OR4 OR4_187 (.A(sel_R_DATA_TEMPR48[19] ), .B(sel_R_DATA_TEMPR49[19] ), 
        .C(sel_R_DATA_TEMPR50[19] ), .D(sel_R_DATA_TEMPR51[19] ), .Y(
        OR4_187_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%51%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R51C0 (.A_DOUT({
        nc152, nc153, nc154, nc155, nc156,int_R_DATA_TEMPR51[31] , 
       int_R_DATA_TEMPR51[30] ,int_R_DATA_TEMPR51[29] , 
       int_R_DATA_TEMPR51[28] ,int_R_DATA_TEMPR51[27] , 
       int_R_DATA_TEMPR51[26] ,int_R_DATA_TEMPR51[25] , 
       int_R_DATA_TEMPR51[24] ,int_R_DATA_TEMPR51[23] , 
       int_R_DATA_TEMPR51[22] ,int_R_DATA_TEMPR51[21] , 
       int_R_DATA_TEMPR51[20] ,int_R_DATA_TEMPR51[19] , 
       int_R_DATA_TEMPR51[18] ,int_R_DATA_TEMPR51[17] }), .B_DOUT({nc157, 
        nc158, nc159,int_R_DATA_TEMPR51[16] ,int_R_DATA_TEMPR51[15] , 
       int_R_DATA_TEMPR51[14] ,int_R_DATA_TEMPR51[13] , 
       int_R_DATA_TEMPR51[12] ,int_R_DATA_TEMPR51[11] , 
       int_R_DATA_TEMPR51[10] ,int_R_DATA_TEMPR51[9] ,int_R_DATA_TEMPR51[8] , 
       int_R_DATA_TEMPR51[7] ,int_R_DATA_TEMPR51[6] ,int_R_DATA_TEMPR51[5] , 
       int_R_DATA_TEMPR51[4] ,int_R_DATA_TEMPR51[3] ,int_R_DATA_TEMPR51[2] , 
       int_R_DATA_TEMPR51[1] ,int_R_DATA_TEMPR51[0] }), .DB_DETECT( int_DB_DETECT_NG[51] ), .SB_CORRECT(int_SB_CORRECT_NG[51] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[51] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[12] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[12] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%79%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R79C0 (.A_DOUT({
        nc160, nc161, nc162, nc163, nc164,int_R_DATA_TEMPR79[31] , 
       int_R_DATA_TEMPR79[30] ,int_R_DATA_TEMPR79[29] , 
       int_R_DATA_TEMPR79[28] ,int_R_DATA_TEMPR79[27] , 
       int_R_DATA_TEMPR79[26] ,int_R_DATA_TEMPR79[25] , 
       int_R_DATA_TEMPR79[24] ,int_R_DATA_TEMPR79[23] , 
       int_R_DATA_TEMPR79[22] ,int_R_DATA_TEMPR79[21] , 
       int_R_DATA_TEMPR79[20] ,int_R_DATA_TEMPR79[19] , 
       int_R_DATA_TEMPR79[18] ,int_R_DATA_TEMPR79[17] }), .B_DOUT({nc165, 
        nc166, nc167,int_R_DATA_TEMPR79[16] ,int_R_DATA_TEMPR79[15] , 
       int_R_DATA_TEMPR79[14] ,int_R_DATA_TEMPR79[13] , 
       int_R_DATA_TEMPR79[12] ,int_R_DATA_TEMPR79[11] , 
       int_R_DATA_TEMPR79[10] ,int_R_DATA_TEMPR79[9] ,int_R_DATA_TEMPR79[8] , 
       int_R_DATA_TEMPR79[7] ,int_R_DATA_TEMPR79[6] ,int_R_DATA_TEMPR79[5] , 
       int_R_DATA_TEMPR79[4] ,int_R_DATA_TEMPR79[3] ,int_R_DATA_TEMPR79[2] , 
       int_R_DATA_TEMPR79[1] ,int_R_DATA_TEMPR79[0] }), .DB_DETECT( int_DB_DETECT_NG[79] ), .SB_CORRECT(int_SB_CORRECT_NG[79] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[79] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[19] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[19] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1052 (.A(OR4_456_Y), .B(OR4_657_Y), .C(OR4_246_Y), .D(
        OR4_19_Y), .Y(OR4_1052_Y));
    OR4 OR4_212 (.A(sel_R_DATA_TEMPR28[7] ), .B(sel_R_DATA_TEMPR29[7] ), .C(sel_R_DATA_TEMPR30[7] ), .D(sel_R_DATA_TEMPR31[7] ), .Y(OR4_212_Y));
    OR4 OR4_1197 (.A(OR4_573_Y), .B(OR4_450_Y), .C(OR4_546_Y), .D(
        OR4_631_Y), .Y(OR4_1197_Y));
    OR4 OR4_353 (.A(OR4_721_Y), .B(OR2_27_Y), .C(sel_R_DATA_TEMPR86[6] ), 
        .D(sel_R_DATA_TEMPR87[6] ), .Y(OR4_353_Y));
    OR4 OR4_1139 (.A(\DB_DETECT[52] ), .B(\DB_DETECT[53] ), .C(
        \DB_DETECT[54] ), .D(\DB_DETECT[55] ), .Y(OR4_1139_Y));
    OR4 OR4_750 (.A(sel_R_DATA_TEMPR120[16] ), .B(sel_R_DATA_TEMPR121[16] ), 
        .C(sel_R_DATA_TEMPR122[16] ), .D(sel_R_DATA_TEMPR123[16] ), .Y(
        OR4_750_Y));
    OR4 OR4_1260 (.A(OR4_695_Y), .B(OR4_556_Y), .C(OR4_49_Y), .D(
        OR4_491_Y), .Y(OR4_1260_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[2]  (.A(CFG3_0_Y), .B(CFG3_2_Y), 
        .Y(\BLKY2[2] ));
    OR4 OR4_783 (.A(sel_R_DATA_TEMPR56[27] ), .B(sel_R_DATA_TEMPR57[27] ), 
        .C(sel_R_DATA_TEMPR58[27] ), .D(sel_R_DATA_TEMPR59[27] ), .Y(
        OR4_783_Y));
    AND4 \AND4SB_CORRECT[90]  (.A(sel_SB_CORRECT_NG[90] ), .B(
        \BLKY2_pipe[22] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[90] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%121%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R121C0 (.A_DOUT({
        nc168, nc169, nc170, nc171, nc172,int_R_DATA_TEMPR121[31] , 
       int_R_DATA_TEMPR121[30] ,int_R_DATA_TEMPR121[29] , 
       int_R_DATA_TEMPR121[28] ,int_R_DATA_TEMPR121[27] , 
       int_R_DATA_TEMPR121[26] ,int_R_DATA_TEMPR121[25] , 
       int_R_DATA_TEMPR121[24] ,int_R_DATA_TEMPR121[23] , 
       int_R_DATA_TEMPR121[22] ,int_R_DATA_TEMPR121[21] , 
       int_R_DATA_TEMPR121[20] ,int_R_DATA_TEMPR121[19] , 
       int_R_DATA_TEMPR121[18] ,int_R_DATA_TEMPR121[17] }), .B_DOUT({nc173, 
        nc174, nc175,int_R_DATA_TEMPR121[16] ,int_R_DATA_TEMPR121[15] , 
       int_R_DATA_TEMPR121[14] ,int_R_DATA_TEMPR121[13] , 
       int_R_DATA_TEMPR121[12] ,int_R_DATA_TEMPR121[11] , 
       int_R_DATA_TEMPR121[10] ,int_R_DATA_TEMPR121[9] , 
       int_R_DATA_TEMPR121[8] ,int_R_DATA_TEMPR121[7] , 
       int_R_DATA_TEMPR121[6] ,int_R_DATA_TEMPR121[5] , 
       int_R_DATA_TEMPR121[4] ,int_R_DATA_TEMPR121[3] , 
       int_R_DATA_TEMPR121[2] ,int_R_DATA_TEMPR121[1] , 
       int_R_DATA_TEMPR121[0] }), .DB_DETECT(int_DB_DETECT_NG[121] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[121] ), .ACCESS_BUSY(
        ACCESS_BUSY[121] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[30] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[30] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1276 (.A(OR4_396_Y), .B(OR4_768_Y), .C(OR4_214_Y), .D(
        OR4_478_Y), .Y(OR4_1276_Y));
    OR4 OR4_600 (.A(sel_R_DATA_TEMPR72[18] ), .B(sel_R_DATA_TEMPR73[18] ), 
        .C(sel_R_DATA_TEMPR74[18] ), .D(sel_R_DATA_TEMPR75[18] ), .Y(
        OR4_600_Y));
    AND4 \AND4DB_DETECT[118]  (.A(sel_DB_DETECT_NG[118] ), .B(
        \BLKY2_pipe[29] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[118] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%37%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R37C0 (.A_DOUT({
        nc176, nc177, nc178, nc179, nc180,int_R_DATA_TEMPR37[31] , 
       int_R_DATA_TEMPR37[30] ,int_R_DATA_TEMPR37[29] , 
       int_R_DATA_TEMPR37[28] ,int_R_DATA_TEMPR37[27] , 
       int_R_DATA_TEMPR37[26] ,int_R_DATA_TEMPR37[25] , 
       int_R_DATA_TEMPR37[24] ,int_R_DATA_TEMPR37[23] , 
       int_R_DATA_TEMPR37[22] ,int_R_DATA_TEMPR37[21] , 
       int_R_DATA_TEMPR37[20] ,int_R_DATA_TEMPR37[19] , 
       int_R_DATA_TEMPR37[18] ,int_R_DATA_TEMPR37[17] }), .B_DOUT({nc181, 
        nc182, nc183,int_R_DATA_TEMPR37[16] ,int_R_DATA_TEMPR37[15] , 
       int_R_DATA_TEMPR37[14] ,int_R_DATA_TEMPR37[13] , 
       int_R_DATA_TEMPR37[12] ,int_R_DATA_TEMPR37[11] , 
       int_R_DATA_TEMPR37[10] ,int_R_DATA_TEMPR37[9] ,int_R_DATA_TEMPR37[8] , 
       int_R_DATA_TEMPR37[7] ,int_R_DATA_TEMPR37[6] ,int_R_DATA_TEMPR37[5] , 
       int_R_DATA_TEMPR37[4] ,int_R_DATA_TEMPR37[3] ,int_R_DATA_TEMPR37[2] , 
       int_R_DATA_TEMPR37[1] ,int_R_DATA_TEMPR37[0] }), .DB_DETECT( int_DB_DETECT_NG[37] ), .SB_CORRECT(int_SB_CORRECT_NG[37] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[37] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[9] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_452 (.A(OR4_641_Y), .B(OR4_903_Y), .C(OR4_1119_Y), .D(
        OR4_944_Y), .Y(OR4_452_Y));
    OR4 OR4_284 (.A(OR4_807_Y), .B(OR4_1073_Y), .C(OR4_603_Y), .D(
        OR4_1341_Y), .Y(OR4_284_Y));
    OR4 OR4_310 (.A(sel_R_DATA_TEMPR64[25] ), .B(sel_R_DATA_TEMPR65[25] ), 
        .C(sel_R_DATA_TEMPR66[25] ), .D(sel_R_DATA_TEMPR67[25] ), .Y(
        OR4_310_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[20]  (.D(\BLKY2[20] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[20] ));
    OR4 OR4_5 (.A(sel_R_DATA_TEMPR16[1] ), .B(sel_R_DATA_TEMPR17[1] ), .C(sel_R_DATA_TEMPR18[1] ), .D(sel_R_DATA_TEMPR19[1] ), .Y(OR4_5_Y));
    OR4 OR4_1316 (.A(OR4_1089_Y), .B(OR4_1393_Y), .C(OR4_145_Y), .D(
        OR4_1166_Y), .Y(OR4_1316_Y));
    AND4 \AND4DB_DETECT[20]  (.A(sel_DB_DETECT_NG[20] ), .B(
        \BLKY2_pipe[5] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[20] ));
    OR4 OR4_1378 (.A(sel_R_DATA_TEMPR56[28] ), .B(sel_R_DATA_TEMPR57[28] ), 
        .C(sel_R_DATA_TEMPR58[28] ), .D(sel_R_DATA_TEMPR59[28] ), .Y(
        OR4_1378_Y));
    OR4 OR4_1046 (.A(OR4_853_Y), .B(OR4_1083_Y), .C(OR4_1259_Y), .D(
        OR4_716_Y), .Y(OR4_1046_Y));
    OR4 OR4_670 (.A(OR4_182_Y), .B(OR2_33_Y), .C(sel_R_DATA_TEMPR86[31] ), 
        .D(sel_R_DATA_TEMPR87[31] ), .Y(OR4_670_Y));
    OR4 OR4_459 (.A(sel_R_DATA_TEMPR40[23] ), .B(sel_R_DATA_TEMPR41[23] ), 
        .C(sel_R_DATA_TEMPR42[23] ), .D(sel_R_DATA_TEMPR43[23] ), .Y(
        OR4_459_Y));
    AND4 \AND4SB_CORRECT[39]  (.A(sel_SB_CORRECT_NG[39] ), .B(
        \BLKY2_pipe[9] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[39] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[27]  (.A(CFG3_19_Y), .B(
        CFG3_3_Y), .Y(\BLKY2[27] ));
    OR4 OR4_307 (.A(sel_R_DATA_TEMPR124[4] ), .B(sel_R_DATA_TEMPR125[4] ), 
        .C(sel_R_DATA_TEMPR126[4] ), .D(sel_R_DATA_TEMPR127[4] ), .Y(
        OR4_307_Y));
    OR4 OR4_100 (.A(OR4_264_Y), .B(OR4_1139_Y), .C(OR4_420_Y), .D(
        OR4_1292_Y), .Y(OR4_100_Y));
    OR4 OR4_1362 (.A(sel_R_DATA_TEMPR96[15] ), .B(sel_R_DATA_TEMPR97[15] ), 
        .C(sel_R_DATA_TEMPR98[15] ), .D(sel_R_DATA_TEMPR99[15] ), .Y(
        OR4_1362_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[28]  (.A(CFG3_6_Y), .B(CFG3_7_Y)
        , .Y(\BLKX2[28] ));
    OR4 OR4_99 (.A(sel_R_DATA_TEMPR104[31] ), .B(sel_R_DATA_TEMPR105[31] ), 
        .C(sel_R_DATA_TEMPR106[31] ), .D(sel_R_DATA_TEMPR107[31] ), .Y(
        OR4_99_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%92%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R92C0 (.A_DOUT({
        nc184, nc185, nc186, nc187, nc188,int_R_DATA_TEMPR92[31] , 
       int_R_DATA_TEMPR92[30] ,int_R_DATA_TEMPR92[29] , 
       int_R_DATA_TEMPR92[28] ,int_R_DATA_TEMPR92[27] , 
       int_R_DATA_TEMPR92[26] ,int_R_DATA_TEMPR92[25] , 
       int_R_DATA_TEMPR92[24] ,int_R_DATA_TEMPR92[23] , 
       int_R_DATA_TEMPR92[22] ,int_R_DATA_TEMPR92[21] , 
       int_R_DATA_TEMPR92[20] ,int_R_DATA_TEMPR92[19] , 
       int_R_DATA_TEMPR92[18] ,int_R_DATA_TEMPR92[17] }), .B_DOUT({nc189, 
        nc190, nc191,int_R_DATA_TEMPR92[16] ,int_R_DATA_TEMPR92[15] , 
       int_R_DATA_TEMPR92[14] ,int_R_DATA_TEMPR92[13] , 
       int_R_DATA_TEMPR92[12] ,int_R_DATA_TEMPR92[11] , 
       int_R_DATA_TEMPR92[10] ,int_R_DATA_TEMPR92[9] ,int_R_DATA_TEMPR92[8] , 
       int_R_DATA_TEMPR92[7] ,int_R_DATA_TEMPR92[6] ,int_R_DATA_TEMPR92[5] , 
       int_R_DATA_TEMPR92[4] ,int_R_DATA_TEMPR92[3] ,int_R_DATA_TEMPR92[2] , 
       int_R_DATA_TEMPR92[1] ,int_R_DATA_TEMPR92[0] }), .DB_DETECT( int_DB_DETECT_NG[92] ), .SB_CORRECT(int_SB_CORRECT_NG[92] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[92] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[23] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[23] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_156 (.A(sel_R_DATA_TEMPR88[4] ), .B(sel_R_DATA_TEMPR89[4] ), .C(sel_R_DATA_TEMPR90[4] ), .D(sel_R_DATA_TEMPR91[4] ), .Y(OR4_156_Y));
    OR4 OR4_1223 (.A(OR4_310_Y), .B(OR4_91_Y), .C(OR4_1240_Y), .D(
        OR4_186_Y), .Y(OR4_1223_Y));
    OR4 OR4_535 (.A(sel_R_DATA_TEMPR72[6] ), .B(sel_R_DATA_TEMPR73[6] ), .C(sel_R_DATA_TEMPR74[6] ), .D(sel_R_DATA_TEMPR75[6] ), .Y(OR4_535_Y));
    OR4 OR4_1262 (.A(OR4_57_Y), .B(OR4_712_Y), .C(OR4_1113_Y), .D(
        OR4_1381_Y), .Y(OR4_1262_Y));
    OR4 OR4_813 (.A(sel_R_DATA_TEMPR92[28] ), .B(sel_R_DATA_TEMPR93[28] ), 
        .C(sel_R_DATA_TEMPR94[28] ), .D(sel_R_DATA_TEMPR95[28] ), .Y(
        OR4_813_Y));
    OR2 OR2_24 (.A(sel_R_DATA_TEMPR84[19] ), .B(sel_R_DATA_TEMPR85[19] ), .Y(
        OR2_24_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[23]  (.A(CFG3_23_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[23] ));
    OR4 OR4_68 (.A(sel_R_DATA_TEMPR28[10] ), .B(sel_R_DATA_TEMPR29[10] ), .C(sel_R_DATA_TEMPR30[10] ), .D(sel_R_DATA_TEMPR31[10] ), .Y(OR4_68_Y));
    AND4 \AND4DB_DETECT[46]  (.A(sel_DB_DETECT_NG[46] ), .B(
        \BLKY2_pipe[11] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[46] ));
    OR4 OR4_377 (.A(sel_R_DATA_TEMPR60[17] ), .B(sel_R_DATA_TEMPR61[17] ), 
        .C(sel_R_DATA_TEMPR62[17] ), .D(sel_R_DATA_TEMPR63[17] ), .Y(
        OR4_377_Y));
    OR4 OR4_170 (.A(sel_R_DATA_TEMPR24[30] ), .B(sel_R_DATA_TEMPR25[30] ), 
        .C(sel_R_DATA_TEMPR26[30] ), .D(sel_R_DATA_TEMPR27[30] ), .Y(
        OR4_170_Y));
    OR4 OR4_1341 (.A(sel_R_DATA_TEMPR60[8] ), .B(sel_R_DATA_TEMPR61[8] ), .C(sel_R_DATA_TEMPR62[8] ), .D(sel_R_DATA_TEMPR63[8] ), .Y(OR4_1341_Y));
    OR4 OR4_708 (.A(sel_R_DATA_TEMPR4[17] ), .B(sel_R_DATA_TEMPR5[17] ), .C(sel_R_DATA_TEMPR6[17] ), .D(sel_R_DATA_TEMPR7[17] ), .Y(OR4_708_Y));
    OR4 OR4_626 (.A(sel_R_DATA_TEMPR76[4] ), .B(sel_R_DATA_TEMPR77[4] ), .C(sel_R_DATA_TEMPR78[4] ), .D(sel_R_DATA_TEMPR79[4] ), .Y(OR4_626_Y));
    OR4 OR4_31 (.A(OR4_295_Y), .B(OR4_69_Y), .C(OR4_1222_Y), .D(
        OR4_521_Y), .Y(OR4_31_Y));
    AND4 \AND4DB_DETECT[41]  (.A(sel_DB_DETECT_NG[41] ), .B(
        \BLKY2_pipe[10] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[41] ));
    DFN1E1 \DFN1E1BLKY2_pipe[31]  (.D(\BLKY2[31] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[31] ));
    AND4 \AND4DB_DETECT[1]  (.A(sel_DB_DETECT_NG[1] ), .B(
        \BLKY2_pipe[0] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[1] ));
    OR4 OR4_633 (.A(sel_R_DATA_TEMPR92[20] ), .B(sel_R_DATA_TEMPR93[20] ), 
        .C(sel_R_DATA_TEMPR94[20] ), .D(sel_R_DATA_TEMPR95[20] ), .Y(
        OR4_633_Y));
    OR4 \OR4_R_DATA[31]  (.A(OR4_324_Y), .B(OR4_261_Y), .C(OR4_283_Y), 
        .D(OR4_1245_Y), .Y(R_DATA[31]));
    AND4 \AND4SB_CORRECT[27]  (.A(sel_SB_CORRECT_NG[27] ), .B(
        \BLKY2_pipe[6] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[27] ));
    OR4 OR4_1136 (.A(OR4_971_Y), .B(OR4_472_Y), .C(OR4_667_Y), .D(
        OR4_1170_Y), .Y(OR4_1136_Y));
    OR4 OR4_385 (.A(OR4_1030_Y), .B(OR4_128_Y), .C(OR4_791_Y), .D(
        OR4_1019_Y), .Y(OR4_385_Y));
    OR4 OR4_778 (.A(sel_R_DATA_TEMPR104[8] ), .B(sel_R_DATA_TEMPR105[8] ), 
        .C(sel_R_DATA_TEMPR106[8] ), .D(sel_R_DATA_TEMPR107[8] ), .Y(
        OR4_778_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[15]  (.A(CFG3_23_Y), .B(
        CFG3_4_Y), .Y(\BLKX2[15] ));
    OR4 OR4_243 (.A(OR4_443_Y), .B(OR4_647_Y), .C(OR4_802_Y), .D(
        OR4_1009_Y), .Y(OR4_243_Y));
    OR4 OR4_394 (.A(\SB_CORRECT[80] ), .B(\SB_CORRECT[81] ), .C(
        \SB_CORRECT[82] ), .D(\SB_CORRECT[83] ), .Y(OR4_394_Y));
    OR4 OR4_1079 (.A(OR4_13_Y), .B(OR4_736_Y), .C(OR4_32_Y), .D(
        OR4_260_Y), .Y(OR4_1079_Y));
    OR4 OR4_1264 (.A(sel_R_DATA_TEMPR100[8] ), .B(sel_R_DATA_TEMPR101[8] ), 
        .C(sel_R_DATA_TEMPR102[8] ), .D(sel_R_DATA_TEMPR103[8] ), .Y(
        OR4_1264_Y));
    OR4 OR4_358 (.A(sel_R_DATA_TEMPR96[26] ), .B(sel_R_DATA_TEMPR97[26] ), 
        .C(sel_R_DATA_TEMPR98[26] ), .D(sel_R_DATA_TEMPR99[26] ), .Y(
        OR4_358_Y));
    OR4 OR4_1231 (.A(OR4_1219_Y), .B(OR4_634_Y), .C(OR4_1091_Y), .D(
        OR4_95_Y), .Y(OR4_1231_Y));
    OR4 OR4_1138 (.A(sel_R_DATA_TEMPR48[29] ), .B(sel_R_DATA_TEMPR49[29] ), 
        .C(sel_R_DATA_TEMPR50[29] ), .D(sel_R_DATA_TEMPR51[29] ), .Y(
        OR4_1138_Y));
    OR4 OR4_80 (.A(sel_R_DATA_TEMPR124[17] ), .B(sel_R_DATA_TEMPR125[17] ), 
        .C(sel_R_DATA_TEMPR126[17] ), .D(sel_R_DATA_TEMPR127[17] ), .Y(
        OR4_80_Y));
    OR4 OR4_1367 (.A(sel_R_DATA_TEMPR48[26] ), .B(sel_R_DATA_TEMPR49[26] ), 
        .C(sel_R_DATA_TEMPR50[26] ), .D(sel_R_DATA_TEMPR51[26] ), .Y(
        OR4_1367_Y));
    OR4 OR4_807 (.A(sel_R_DATA_TEMPR48[8] ), .B(sel_R_DATA_TEMPR49[8] ), .C(sel_R_DATA_TEMPR50[8] ), .D(sel_R_DATA_TEMPR51[8] ), .Y(OR4_807_Y));
    OR4 OR4_108 (.A(OR4_611_Y), .B(OR2_31_Y), .C(sel_R_DATA_TEMPR86[12] ), 
        .D(sel_R_DATA_TEMPR87[12] ), .Y(OR4_108_Y));
    OR4 OR4_191 (.A(sel_R_DATA_TEMPR16[12] ), .B(sel_R_DATA_TEMPR17[12] ), 
        .C(sel_R_DATA_TEMPR18[12] ), .D(sel_R_DATA_TEMPR19[12] ), .Y(
        OR4_191_Y));
    OR4 OR4_1290 (.A(sel_R_DATA_TEMPR68[2] ), .B(sel_R_DATA_TEMPR69[2] ), .C(sel_R_DATA_TEMPR70[2] ), .D(sel_R_DATA_TEMPR71[2] ), .Y(OR4_1290_Y));
    OR4 OR4_1129 (.A(OR4_1266_Y), .B(OR4_94_Y), .C(OR4_253_Y), .D(
        OR4_1342_Y), .Y(OR4_1129_Y));
    OR4 OR4_904 (.A(OR4_1365_Y), .B(OR4_185_Y), .C(OR4_1158_Y), .D(
        OR4_928_Y), .Y(OR4_904_Y));
    OR4 OR4_948 (.A(sel_R_DATA_TEMPR124[26] ), .B(sel_R_DATA_TEMPR125[26] ), 
        .C(sel_R_DATA_TEMPR126[26] ), .D(sel_R_DATA_TEMPR127[26] ), .Y(
        OR4_948_Y));
    OR4 OR4_1 (.A(sel_R_DATA_TEMPR44[28] ), .B(sel_R_DATA_TEMPR45[28] ), .C(sel_R_DATA_TEMPR46[28] ), .D(sel_R_DATA_TEMPR47[28] ), .Y(OR4_1_Y));
    AND4 \AND4DB_DETECT[18]  (.A(sel_DB_DETECT_NG[18] ), .B(
        \BLKY2_pipe[4] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[18] ));
    OR4 OR4_87 (.A(sel_R_DATA_TEMPR96[18] ), .B(sel_R_DATA_TEMPR97[18] ), .C(sel_R_DATA_TEMPR98[18] ), .D(sel_R_DATA_TEMPR99[18] ), .Y(OR4_87_Y));
    OR4 OR4_877 (.A(sel_R_DATA_TEMPR116[29] ), .B(sel_R_DATA_TEMPR117[29] ), 
        .C(sel_R_DATA_TEMPR118[29] ), .D(sel_R_DATA_TEMPR119[29] ), .Y(
        OR4_877_Y));
    OR4 \OR4_R_DATA[30]  (.A(OR4_71_Y), .B(OR4_378_Y), .C(OR4_1003_Y), 
        .D(OR4_482_Y), .Y(R_DATA[30]));
    OR4 OR4_178 (.A(sel_R_DATA_TEMPR8[7] ), .B(sel_R_DATA_TEMPR9[7] ), .C(sel_R_DATA_TEMPR10[7] ), .D(sel_R_DATA_TEMPR11[7] ), .Y(OR4_178_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[0]  (.A(CFG3_13_Y), .B(
        CFG3_12_Y), .Y(\BLKX2[0] ));
    OR4 OR4_974 (.A(sel_R_DATA_TEMPR124[13] ), .B(sel_R_DATA_TEMPR125[13] ), 
        .C(sel_R_DATA_TEMPR126[13] ), .D(sel_R_DATA_TEMPR127[13] ), .Y(
        OR4_974_Y));
    OR4 OR4_939 (.A(sel_R_DATA_TEMPR32[14] ), .B(sel_R_DATA_TEMPR33[14] ), 
        .C(sel_R_DATA_TEMPR34[14] ), .D(sel_R_DATA_TEMPR35[14] ), .Y(
        OR4_939_Y));
    OR4 OR4_930 (.A(sel_R_DATA_TEMPR80[21] ), .B(sel_R_DATA_TEMPR81[21] ), 
        .C(sel_R_DATA_TEMPR82[21] ), .D(sel_R_DATA_TEMPR83[21] ), .Y(
        OR4_930_Y));
    AND4 \AND4SB_CORRECT[83]  (.A(sel_SB_CORRECT_NG[83] ), .B(
        \BLKY2_pipe[20] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[83] ));
    AND4 \AND4DB_DETECT[97]  (.A(sel_DB_DETECT_NG[97] ), .B(
        \BLKY2_pipe[24] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[97] ));
    OR4 OR4_1392 (.A(OR4_729_Y), .B(OR4_1192_Y), .C(OR4_303_Y), .D(
        OR4_100_Y), .Y(OR4_1392_Y));
    OR4 OR4_782 (.A(sel_R_DATA_TEMPR64[24] ), .B(sel_R_DATA_TEMPR65[24] ), 
        .C(sel_R_DATA_TEMPR66[24] ), .D(sel_R_DATA_TEMPR67[24] ), .Y(
        OR4_782_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[11]  (.D(\BLKY2[11] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[11] ));
    OR4 OR4_159 (.A(sel_R_DATA_TEMPR64[6] ), .B(sel_R_DATA_TEMPR65[6] ), .C(sel_R_DATA_TEMPR66[6] ), .D(sel_R_DATA_TEMPR67[6] ), .Y(OR4_159_Y));
    OR4 OR4_491 (.A(sel_R_DATA_TEMPR60[31] ), .B(sel_R_DATA_TEMPR61[31] ), 
        .C(sel_R_DATA_TEMPR62[31] ), .D(sel_R_DATA_TEMPR63[31] ), .Y(
        OR4_491_Y));
    OR4 OR4_165 (.A(sel_R_DATA_TEMPR12[6] ), .B(sel_R_DATA_TEMPR13[6] ), .C(sel_R_DATA_TEMPR14[6] ), .D(sel_R_DATA_TEMPR15[6] ), .Y(OR4_165_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%46%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R46C0 (.A_DOUT({
        nc192, nc193, nc194, nc195, nc196,int_R_DATA_TEMPR46[31] , 
       int_R_DATA_TEMPR46[30] ,int_R_DATA_TEMPR46[29] , 
       int_R_DATA_TEMPR46[28] ,int_R_DATA_TEMPR46[27] , 
       int_R_DATA_TEMPR46[26] ,int_R_DATA_TEMPR46[25] , 
       int_R_DATA_TEMPR46[24] ,int_R_DATA_TEMPR46[23] , 
       int_R_DATA_TEMPR46[22] ,int_R_DATA_TEMPR46[21] , 
       int_R_DATA_TEMPR46[20] ,int_R_DATA_TEMPR46[19] , 
       int_R_DATA_TEMPR46[18] ,int_R_DATA_TEMPR46[17] }), .B_DOUT({nc197, 
        nc198, nc199,int_R_DATA_TEMPR46[16] ,int_R_DATA_TEMPR46[15] , 
       int_R_DATA_TEMPR46[14] ,int_R_DATA_TEMPR46[13] , 
       int_R_DATA_TEMPR46[12] ,int_R_DATA_TEMPR46[11] , 
       int_R_DATA_TEMPR46[10] ,int_R_DATA_TEMPR46[9] ,int_R_DATA_TEMPR46[8] , 
       int_R_DATA_TEMPR46[7] ,int_R_DATA_TEMPR46[6] ,int_R_DATA_TEMPR46[5] , 
       int_R_DATA_TEMPR46[4] ,int_R_DATA_TEMPR46[3] ,int_R_DATA_TEMPR46[2] , 
       int_R_DATA_TEMPR46[1] ,int_R_DATA_TEMPR46[0] }), .DB_DETECT( int_DB_DETECT_NG[46] ), .SB_CORRECT(int_SB_CORRECT_NG[46] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[46] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[11] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[11] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1292 (.A(\DB_DETECT[60] ), .B(\DB_DETECT[61] ), .C(
        \DB_DETECT[62] ), .D(\DB_DETECT[63] ), .Y(OR4_1292_Y));
    OR4 OR4_133 (.A(sel_R_DATA_TEMPR120[28] ), .B(sel_R_DATA_TEMPR121[28] ), 
        .C(sel_R_DATA_TEMPR122[28] ), .D(sel_R_DATA_TEMPR123[28] ), .Y(
        OR4_133_Y));
    OR4 OR4_515 (.A(sel_R_DATA_TEMPR40[19] ), .B(sel_R_DATA_TEMPR41[19] ), 
        .C(sel_R_DATA_TEMPR42[19] ), .D(sel_R_DATA_TEMPR43[19] ), .Y(
        OR4_515_Y));
    OR4 OR4_498 (.A(sel_R_DATA_TEMPR96[30] ), .B(sel_R_DATA_TEMPR97[30] ), 
        .C(sel_R_DATA_TEMPR98[30] ), .D(sel_R_DATA_TEMPR99[30] ), .Y(
        OR4_498_Y));
    AND4 \AND4DB_DETECT[67]  (.A(sel_DB_DETECT_NG[67] ), .B(
        \BLKY2_pipe[16] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[67] ));
    OR4 OR4_986 (.A(sel_R_DATA_TEMPR64[7] ), .B(sel_R_DATA_TEMPR65[7] ), .C(sel_R_DATA_TEMPR66[7] ), .D(sel_R_DATA_TEMPR67[7] ), .Y(OR4_986_Y));
    OR4 OR4_467 (.A(OR4_905_Y), .B(OR4_1180_Y), .C(OR4_694_Y), .D(
        OR4_48_Y), .Y(OR4_467_Y));
    AND4 \AND4SB_CORRECT[67]  (.A(sel_SB_CORRECT_NG[67] ), .B(
        \BLKY2_pipe[16] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[67] ));
    OR4 OR4_92 (.A(sel_R_DATA_TEMPR60[15] ), .B(sel_R_DATA_TEMPR61[15] ), .C(sel_R_DATA_TEMPR62[15] ), .D(sel_R_DATA_TEMPR63[15] ), .Y(OR4_92_Y));
    OR4 OR4_1103 (.A(sel_R_DATA_TEMPR52[10] ), .B(sel_R_DATA_TEMPR53[10] ), 
        .C(sel_R_DATA_TEMPR54[10] ), .D(sel_R_DATA_TEMPR55[10] ), .Y(
        OR4_1103_Y));
    OR4 OR4_648 (.A(sel_R_DATA_TEMPR56[19] ), .B(sel_R_DATA_TEMPR57[19] ), 
        .C(sel_R_DATA_TEMPR58[19] ), .D(sel_R_DATA_TEMPR59[19] ), .Y(
        OR4_648_Y));
    OR4 OR4_1114 (.A(sel_R_DATA_TEMPR112[29] ), .B(sel_R_DATA_TEMPR113[29] ), 
        .C(sel_R_DATA_TEMPR114[29] ), .D(sel_R_DATA_TEMPR115[29] ), .Y(
        OR4_1114_Y));
    OR4 OR4_685 (.A(sel_R_DATA_TEMPR68[10] ), .B(sel_R_DATA_TEMPR69[10] ), 
        .C(sel_R_DATA_TEMPR70[10] ), .D(sel_R_DATA_TEMPR71[10] ), .Y(
        OR4_685_Y));
    AND4 \AND4DB_DETECT[109]  (.A(sel_DB_DETECT_NG[109] ), .B(
        \BLKY2_pipe[27] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[109] ));
    AND4 \AND4DB_DETECT[55]  (.A(sel_DB_DETECT_NG[55] ), .B(
        \BLKY2_pipe[13] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[55] ));
    OR4 OR4_613 (.A(OR4_707_Y), .B(OR4_494_Y), .C(OR4_249_Y), .D(
        OR4_744_Y), .Y(OR4_613_Y));
    OR4 OR4_1126 (.A(sel_R_DATA_TEMPR56[26] ), .B(sel_R_DATA_TEMPR57[26] ), 
        .C(sel_R_DATA_TEMPR58[26] ), .D(sel_R_DATA_TEMPR59[26] ), .Y(
        OR4_1126_Y));
    OR4 OR4_951 (.A(OR4_756_Y), .B(OR4_781_Y), .C(OR4_760_Y), .D(
        OR4_50_Y), .Y(OR4_951_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[28]  (.A(CFG3_18_Y), .B(
        CFG3_3_Y), .Y(\BLKY2[28] ));
    OR4 OR4_642 (.A(OR4_1315_Y), .B(OR4_893_Y), .C(OR4_963_Y), .D(
        OR4_1235_Y), .Y(OR4_642_Y));
    OR4 OR4_1294 (.A(sel_R_DATA_TEMPR72[9] ), .B(sel_R_DATA_TEMPR73[9] ), .C(sel_R_DATA_TEMPR74[9] ), .D(sel_R_DATA_TEMPR75[9] ), .Y(OR4_1294_Y));
    OR2 OR2_30 (.A(sel_R_DATA_TEMPR84[23] ), .B(sel_R_DATA_TEMPR85[23] ), .Y(
        OR2_30_Y));
    AND4 \AND4SB_CORRECT[84]  (.A(sel_SB_CORRECT_NG[84] ), .B(
        \BLKY2_pipe[21] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[84] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%7%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R7C0 (.A_DOUT({
        nc200, nc201, nc202, nc203, nc204,int_R_DATA_TEMPR7[31] , 
       int_R_DATA_TEMPR7[30] ,int_R_DATA_TEMPR7[29] ,int_R_DATA_TEMPR7[28] , 
       int_R_DATA_TEMPR7[27] ,int_R_DATA_TEMPR7[26] ,int_R_DATA_TEMPR7[25] , 
       int_R_DATA_TEMPR7[24] ,int_R_DATA_TEMPR7[23] ,int_R_DATA_TEMPR7[22] , 
       int_R_DATA_TEMPR7[21] ,int_R_DATA_TEMPR7[20] ,int_R_DATA_TEMPR7[19] , 
       int_R_DATA_TEMPR7[18] ,int_R_DATA_TEMPR7[17] }), .B_DOUT({nc205, 
        nc206, nc207,int_R_DATA_TEMPR7[16] ,int_R_DATA_TEMPR7[15] , 
       int_R_DATA_TEMPR7[14] ,int_R_DATA_TEMPR7[13] ,int_R_DATA_TEMPR7[12] , 
       int_R_DATA_TEMPR7[11] ,int_R_DATA_TEMPR7[10] ,int_R_DATA_TEMPR7[9] , 
       int_R_DATA_TEMPR7[8] ,int_R_DATA_TEMPR7[7] ,int_R_DATA_TEMPR7[6] , 
       int_R_DATA_TEMPR7[5] ,int_R_DATA_TEMPR7[4] ,int_R_DATA_TEMPR7[3] , 
       int_R_DATA_TEMPR7[2] ,int_R_DATA_TEMPR7[1] ,int_R_DATA_TEMPR7[0] }), 
        .DB_DETECT(int_DB_DETECT_NG[7] ), .SB_CORRECT( int_SB_CORRECT_NG[7] ), .ACCESS_BUSY(\ACCESS_BUSY[7] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[1] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1221 (.A(sel_R_DATA_TEMPR116[15] ), .B(sel_R_DATA_TEMPR117[15] ), 
        .C(sel_R_DATA_TEMPR118[15] ), .D(sel_R_DATA_TEMPR119[15] ), .Y(
        OR4_1221_Y));
    OR4 OR4_324 (.A(OR4_779_Y), .B(OR4_1023_Y), .C(OR4_1018_Y), .D(
        OR4_1260_Y), .Y(OR4_324_Y));
    OR4 OR4_265 (.A(OR4_56_Y), .B(OR4_1228_Y), .C(OR4_961_Y), .D(
        OR4_1088_Y), .Y(OR4_265_Y));
    OR4 OR4_1128 (.A(sel_R_DATA_TEMPR68[9] ), .B(sel_R_DATA_TEMPR69[9] ), .C(sel_R_DATA_TEMPR70[9] ), .D(sel_R_DATA_TEMPR71[9] ), .Y(OR4_1128_Y));
    OR4 OR4_49 (.A(sel_R_DATA_TEMPR56[31] ), .B(sel_R_DATA_TEMPR57[31] ), .C(sel_R_DATA_TEMPR58[31] ), .D(sel_R_DATA_TEMPR59[31] ), .Y(OR4_49_Y));
    OR4 OR4_599 (.A(OR4_628_Y), .B(OR4_886_Y), .C(OR4_434_Y), .D(
        OR4_1155_Y), .Y(OR4_599_Y));
    OR2 OR2_14 (.A(sel_R_DATA_TEMPR84[8] ), .B(sel_R_DATA_TEMPR85[8] ), .Y(
        OR2_14_Y));
    OR4 OR4_1218 (.A(OR4_364_Y), .B(OR4_1171_Y), .C(OR4_1241_Y), .D(
        OR4_543_Y), .Y(OR4_1218_Y));
    OR4 OR4_862 (.A(OR4_703_Y), .B(OR2_6_Y), .C(sel_R_DATA_TEMPR86[28] ), 
        .D(sel_R_DATA_TEMPR87[28] ), .Y(OR4_862_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[23]  (.A(CFG3_21_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[23] ));
    OR4 OR4_590 (.A(sel_R_DATA_TEMPR28[4] ), .B(sel_R_DATA_TEMPR29[4] ), .C(sel_R_DATA_TEMPR30[4] ), .D(sel_R_DATA_TEMPR31[4] ), .Y(OR4_590_Y));
    OR4 OR4_121 (.A(sel_R_DATA_TEMPR80[8] ), .B(sel_R_DATA_TEMPR81[8] ), .C(sel_R_DATA_TEMPR82[8] ), .D(sel_R_DATA_TEMPR83[8] ), .Y(OR4_121_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[5]  (.A(CFG3_22_Y), .B(
        CFG3_12_Y), .Y(\BLKX2[5] ));
    OR4 OR4_1183 (.A(OR4_231_Y), .B(OR2_18_Y), .C(sel_R_DATA_TEMPR86[0] ), 
        .D(sel_R_DATA_TEMPR87[0] ), .Y(OR4_1183_Y));
    OR4 OR4_1142 (.A(OR4_1090_Y), .B(OR4_1079_Y), .C(OR4_990_Y), .D(
        OR4_1345_Y), .Y(OR4_1142_Y));
    AND4 \AND4DB_DETECT[119]  (.A(sel_DB_DETECT_NG[119] ), .B(
        \BLKY2_pipe[29] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[119] ));
    OR4 OR4_919 (.A(OR4_273_Y), .B(OR4_257_Y), .C(OR4_701_Y), .D(
        OR4_193_Y), .Y(OR4_919_Y));
    OR4 OR4_910 (.A(OR4_620_Y), .B(OR4_833_Y), .C(OR4_996_Y), .D(
        OR4_1057_Y), .Y(OR4_910_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%19%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R19C0 (.A_DOUT({
        nc208, nc209, nc210, nc211, nc212,int_R_DATA_TEMPR19[31] , 
       int_R_DATA_TEMPR19[30] ,int_R_DATA_TEMPR19[29] , 
       int_R_DATA_TEMPR19[28] ,int_R_DATA_TEMPR19[27] , 
       int_R_DATA_TEMPR19[26] ,int_R_DATA_TEMPR19[25] , 
       int_R_DATA_TEMPR19[24] ,int_R_DATA_TEMPR19[23] , 
       int_R_DATA_TEMPR19[22] ,int_R_DATA_TEMPR19[21] , 
       int_R_DATA_TEMPR19[20] ,int_R_DATA_TEMPR19[19] , 
       int_R_DATA_TEMPR19[18] ,int_R_DATA_TEMPR19[17] }), .B_DOUT({nc213, 
        nc214, nc215,int_R_DATA_TEMPR19[16] ,int_R_DATA_TEMPR19[15] , 
       int_R_DATA_TEMPR19[14] ,int_R_DATA_TEMPR19[13] , 
       int_R_DATA_TEMPR19[12] ,int_R_DATA_TEMPR19[11] , 
       int_R_DATA_TEMPR19[10] ,int_R_DATA_TEMPR19[9] ,int_R_DATA_TEMPR19[8] , 
       int_R_DATA_TEMPR19[7] ,int_R_DATA_TEMPR19[6] ,int_R_DATA_TEMPR19[5] , 
       int_R_DATA_TEMPR19[4] ,int_R_DATA_TEMPR19[3] ,int_R_DATA_TEMPR19[2] , 
       int_R_DATA_TEMPR19[1] ,int_R_DATA_TEMPR19[0] }), .DB_DETECT( int_DB_DETECT_NG[19] ), .SB_CORRECT(int_SB_CORRECT_NG[19] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[19] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[4] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 \OR4_R_DATA[18]  (.A(OR4_1320_Y), .B(OR4_1132_Y), .C(OR4_503_Y)
        , .D(OR4_684_Y), .Y(R_DATA[18]));
    AND4 \AND4SB_CORRECT[119]  (.A(sel_SB_CORRECT_NG[119] ), .B(
        \BLKY2_pipe[29] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[119] ));
    OR4 OR4_830 (.A(sel_R_DATA_TEMPR52[13] ), .B(sel_R_DATA_TEMPR53[13] ), 
        .C(sel_R_DATA_TEMPR54[13] ), .D(sel_R_DATA_TEMPR55[13] ), .Y(
        OR4_830_Y));
    OR4 OR4_1177 (.A(OR4_188_Y), .B(OR4_23_Y), .C(OR4_1104_Y), .D(
        OR4_953_Y), .Y(OR4_1177_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%77%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R77C0 (.A_DOUT({
        nc216, nc217, nc218, nc219, nc220,int_R_DATA_TEMPR77[31] , 
       int_R_DATA_TEMPR77[30] ,int_R_DATA_TEMPR77[29] , 
       int_R_DATA_TEMPR77[28] ,int_R_DATA_TEMPR77[27] , 
       int_R_DATA_TEMPR77[26] ,int_R_DATA_TEMPR77[25] , 
       int_R_DATA_TEMPR77[24] ,int_R_DATA_TEMPR77[23] , 
       int_R_DATA_TEMPR77[22] ,int_R_DATA_TEMPR77[21] , 
       int_R_DATA_TEMPR77[20] ,int_R_DATA_TEMPR77[19] , 
       int_R_DATA_TEMPR77[18] ,int_R_DATA_TEMPR77[17] }), .B_DOUT({nc221, 
        nc222, nc223,int_R_DATA_TEMPR77[16] ,int_R_DATA_TEMPR77[15] , 
       int_R_DATA_TEMPR77[14] ,int_R_DATA_TEMPR77[13] , 
       int_R_DATA_TEMPR77[12] ,int_R_DATA_TEMPR77[11] , 
       int_R_DATA_TEMPR77[10] ,int_R_DATA_TEMPR77[9] ,int_R_DATA_TEMPR77[8] , 
       int_R_DATA_TEMPR77[7] ,int_R_DATA_TEMPR77[6] ,int_R_DATA_TEMPR77[5] , 
       int_R_DATA_TEMPR77[4] ,int_R_DATA_TEMPR77[3] ,int_R_DATA_TEMPR77[2] , 
       int_R_DATA_TEMPR77[1] ,int_R_DATA_TEMPR77[0] }), .DB_DETECT( int_DB_DETECT_NG[77] ), .SB_CORRECT(int_SB_CORRECT_NG[77] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[77] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[19] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_680 (.A(sel_R_DATA_TEMPR32[25] ), .B(sel_R_DATA_TEMPR33[25] ), 
        .C(sel_R_DATA_TEMPR34[25] ), .D(sel_R_DATA_TEMPR35[25] ), .Y(
        OR4_680_Y));
    OR4 OR4_113 (.A(OR4_83_Y), .B(OR4_341_Y), .C(OR4_544_Y), .D(
        OR4_384_Y), .Y(OR4_113_Y));
    OR4 OR4_132 (.A(sel_R_DATA_TEMPR28[19] ), .B(sel_R_DATA_TEMPR29[19] ), 
        .C(sel_R_DATA_TEMPR30[19] ), .D(sel_R_DATA_TEMPR31[19] ), .Y(
        OR4_132_Y));
    OR4 OR4_7 (.A(OR4_1029_Y), .B(OR4_126_Y), .C(OR4_790_Y), .D(
        OR4_1017_Y), .Y(OR4_7_Y));
    OR4 OR4_845 (.A(OR4_910_Y), .B(OR4_718_Y), .C(OR4_1186_Y), .D(
        OR4_173_Y), .Y(OR4_845_Y));
    OR4 OR4_421 (.A(OR4_1194_Y), .B(OR4_63_Y), .C(OR4_969_Y), .D(
        OR4_316_Y), .Y(OR4_421_Y));
    OR4 OR4_935 (.A(sel_R_DATA_TEMPR72[4] ), .B(sel_R_DATA_TEMPR73[4] ), .C(sel_R_DATA_TEMPR74[4] ), .D(sel_R_DATA_TEMPR75[4] ), .Y(OR4_935_Y));
    OR4 OR4_463 (.A(sel_R_DATA_TEMPR108[11] ), .B(sel_R_DATA_TEMPR109[11] ), 
        .C(sel_R_DATA_TEMPR110[11] ), .D(sel_R_DATA_TEMPR111[11] ), .Y(
        OR4_463_Y));
    OR4 OR4_755 (.A(sel_R_DATA_TEMPR76[1] ), .B(sel_R_DATA_TEMPR77[1] ), .C(sel_R_DATA_TEMPR78[1] ), .D(sel_R_DATA_TEMPR79[1] ), .Y(OR4_755_Y));
    OR4 OR4_661 (.A(sel_R_DATA_TEMPR52[16] ), .B(sel_R_DATA_TEMPR53[16] ), 
        .C(sel_R_DATA_TEMPR54[16] ), .D(sel_R_DATA_TEMPR55[16] ), .Y(
        OR4_661_Y));
    OR4 OR4_657 (.A(sel_R_DATA_TEMPR20[27] ), .B(sel_R_DATA_TEMPR21[27] ), 
        .C(sel_R_DATA_TEMPR22[27] ), .D(sel_R_DATA_TEMPR23[27] ), .Y(
        OR4_657_Y));
    OR4 OR4_428 (.A(sel_R_DATA_TEMPR12[16] ), .B(sel_R_DATA_TEMPR13[16] ), 
        .C(sel_R_DATA_TEMPR14[16] ), .D(sel_R_DATA_TEMPR15[16] ), .Y(
        OR4_428_Y));
    AND4 \AND4DB_DETECT[102]  (.A(sel_DB_DETECT_NG[102] ), .B(
        \BLKY2_pipe[25] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[102] ));
    AND4 \AND4DB_DETECT[74]  (.A(sel_DB_DETECT_NG[74] ), .B(
        \BLKY2_pipe[18] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[74] ));
    OR4 OR4_1366 (.A(sel_R_DATA_TEMPR40[0] ), .B(sel_R_DATA_TEMPR41[0] ), .C(sel_R_DATA_TEMPR42[0] ), .D(sel_R_DATA_TEMPR43[0] ), .Y(OR4_1366_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%84%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R84C0 (.A_DOUT({
        nc224, nc225, nc226, nc227, nc228,int_R_DATA_TEMPR84[31] , 
       int_R_DATA_TEMPR84[30] ,int_R_DATA_TEMPR84[29] , 
       int_R_DATA_TEMPR84[28] ,int_R_DATA_TEMPR84[27] , 
       int_R_DATA_TEMPR84[26] ,int_R_DATA_TEMPR84[25] , 
       int_R_DATA_TEMPR84[24] ,int_R_DATA_TEMPR84[23] , 
       int_R_DATA_TEMPR84[22] ,int_R_DATA_TEMPR84[21] , 
       int_R_DATA_TEMPR84[20] ,int_R_DATA_TEMPR84[19] , 
       int_R_DATA_TEMPR84[18] ,int_R_DATA_TEMPR84[17] }), .B_DOUT({nc229, 
        nc230, nc231,int_R_DATA_TEMPR84[16] ,int_R_DATA_TEMPR84[15] , 
       int_R_DATA_TEMPR84[14] ,int_R_DATA_TEMPR84[13] , 
       int_R_DATA_TEMPR84[12] ,int_R_DATA_TEMPR84[11] , 
       int_R_DATA_TEMPR84[10] ,int_R_DATA_TEMPR84[9] ,int_R_DATA_TEMPR84[8] , 
       int_R_DATA_TEMPR84[7] ,int_R_DATA_TEMPR84[6] ,int_R_DATA_TEMPR84[5] , 
       int_R_DATA_TEMPR84[4] ,int_R_DATA_TEMPR84[3] ,int_R_DATA_TEMPR84[2] , 
       int_R_DATA_TEMPR84[1] ,int_R_DATA_TEMPR84[0] }), .DB_DETECT( int_DB_DETECT_NG[84] ), .SB_CORRECT(int_SB_CORRECT_NG[84] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[84] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[21] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[21] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4DB_DETECT[28]  (.A(sel_DB_DETECT_NG[28] ), .B(
        \BLKY2_pipe[7] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[28] ));
    OR4 OR4_756 (.A(OR4_74_Y), .B(OR4_1313_Y), .C(OR4_35_Y), .D(
        OR4_550_Y), .Y(OR4_756_Y));
    OR4 OR4_268 (.A(OR4_1352_Y), .B(OR4_62_Y), .C(OR4_517_Y), .D(
        OR4_1_Y), .Y(OR4_268_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%93%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R93C0 (.A_DOUT({
        nc232, nc233, nc234, nc235, nc236,int_R_DATA_TEMPR93[31] , 
       int_R_DATA_TEMPR93[30] ,int_R_DATA_TEMPR93[29] , 
       int_R_DATA_TEMPR93[28] ,int_R_DATA_TEMPR93[27] , 
       int_R_DATA_TEMPR93[26] ,int_R_DATA_TEMPR93[25] , 
       int_R_DATA_TEMPR93[24] ,int_R_DATA_TEMPR93[23] , 
       int_R_DATA_TEMPR93[22] ,int_R_DATA_TEMPR93[21] , 
       int_R_DATA_TEMPR93[20] ,int_R_DATA_TEMPR93[19] , 
       int_R_DATA_TEMPR93[18] ,int_R_DATA_TEMPR93[17] }), .B_DOUT({nc237, 
        nc238, nc239,int_R_DATA_TEMPR93[16] ,int_R_DATA_TEMPR93[15] , 
       int_R_DATA_TEMPR93[14] ,int_R_DATA_TEMPR93[13] , 
       int_R_DATA_TEMPR93[12] ,int_R_DATA_TEMPR93[11] , 
       int_R_DATA_TEMPR93[10] ,int_R_DATA_TEMPR93[9] ,int_R_DATA_TEMPR93[8] , 
       int_R_DATA_TEMPR93[7] ,int_R_DATA_TEMPR93[6] ,int_R_DATA_TEMPR93[5] , 
       int_R_DATA_TEMPR93[4] ,int_R_DATA_TEMPR93[3] ,int_R_DATA_TEMPR93[2] , 
       int_R_DATA_TEMPR93[1] ,int_R_DATA_TEMPR93[0] }), .DB_DETECT( int_DB_DETECT_NG[93] ), .SB_CORRECT(int_SB_CORRECT_NG[93] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[93] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[23] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[23] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_387 (.A(sel_R_DATA_TEMPR108[18] ), .B(sel_R_DATA_TEMPR109[18] ), 
        .C(sel_R_DATA_TEMPR110[18] ), .D(sel_R_DATA_TEMPR111[18] ), .Y(
        OR4_387_Y));
    OR4 OR4_180 (.A(\DB_DETECT[40] ), .B(\DB_DETECT[41] ), .C(
        \DB_DETECT[42] ), .D(\DB_DETECT[43] ), .Y(OR4_180_Y));
    OR4 OR4_105 (.A(OR4_555_Y), .B(OR4_766_Y), .C(OR4_935_Y), .D(
        OR4_626_Y), .Y(OR4_105_Y));
    AND4 \AND4SB_CORRECT[126]  (.A(sel_SB_CORRECT_NG[126] ), .B(
        \BLKY2_pipe[31] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[126] ));
    AND4 \AND4DB_DETECT[19]  (.A(sel_DB_DETECT_NG[19] ), .B(
        \BLKY2_pipe[4] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[19] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%36%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R36C0 (.A_DOUT({
        nc240, nc241, nc242, nc243, nc244,int_R_DATA_TEMPR36[31] , 
       int_R_DATA_TEMPR36[30] ,int_R_DATA_TEMPR36[29] , 
       int_R_DATA_TEMPR36[28] ,int_R_DATA_TEMPR36[27] , 
       int_R_DATA_TEMPR36[26] ,int_R_DATA_TEMPR36[25] , 
       int_R_DATA_TEMPR36[24] ,int_R_DATA_TEMPR36[23] , 
       int_R_DATA_TEMPR36[22] ,int_R_DATA_TEMPR36[21] , 
       int_R_DATA_TEMPR36[20] ,int_R_DATA_TEMPR36[19] , 
       int_R_DATA_TEMPR36[18] ,int_R_DATA_TEMPR36[17] }), .B_DOUT({nc245, 
        nc246, nc247,int_R_DATA_TEMPR36[16] ,int_R_DATA_TEMPR36[15] , 
       int_R_DATA_TEMPR36[14] ,int_R_DATA_TEMPR36[13] , 
       int_R_DATA_TEMPR36[12] ,int_R_DATA_TEMPR36[11] , 
       int_R_DATA_TEMPR36[10] ,int_R_DATA_TEMPR36[9] ,int_R_DATA_TEMPR36[8] , 
       int_R_DATA_TEMPR36[7] ,int_R_DATA_TEMPR36[6] ,int_R_DATA_TEMPR36[5] , 
       int_R_DATA_TEMPR36[4] ,int_R_DATA_TEMPR36[3] ,int_R_DATA_TEMPR36[2] , 
       int_R_DATA_TEMPR36[1] ,int_R_DATA_TEMPR36[0] }), .DB_DETECT( int_DB_DETECT_NG[36] ), .SB_CORRECT(int_SB_CORRECT_NG[36] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[36] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[9] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[9] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_788 (.A(sel_R_DATA_TEMPR4[5] ), .B(sel_R_DATA_TEMPR5[5] ), .C(sel_R_DATA_TEMPR6[5] ), .D(sel_R_DATA_TEMPR7[5] ), .Y(OR4_788_Y));
    OR4 OR4_407 (.A(sel_R_DATA_TEMPR88[30] ), .B(sel_R_DATA_TEMPR89[30] ), 
        .C(sel_R_DATA_TEMPR90[30] ), .D(sel_R_DATA_TEMPR91[30] ), .Y(
        OR4_407_Y));
    AND4 \AND4SB_CORRECT[123]  (.A(sel_SB_CORRECT_NG[123] ), .B(
        \BLKY2_pipe[30] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[123] ));
    CFG3 #( .INIT(8'h10) )  CFG3_15 (.A(R_ADDR[13]), .B(R_ADDR[12]), 
        .C(R_ADDR[11]), .Y(CFG3_15_Y));
    OR4 OR4_175 (.A(sel_R_DATA_TEMPR56[20] ), .B(sel_R_DATA_TEMPR57[20] ), 
        .C(sel_R_DATA_TEMPR58[20] ), .D(sel_R_DATA_TEMPR59[20] ), .Y(
        OR4_175_Y));
    OR4 OR4_393 (.A(sel_R_DATA_TEMPR124[24] ), .B(sel_R_DATA_TEMPR125[24] ), 
        .C(sel_R_DATA_TEMPR126[24] ), .D(sel_R_DATA_TEMPR127[24] ), .Y(
        OR4_393_Y));
    OR4 OR4_790 (.A(sel_R_DATA_TEMPR104[24] ), .B(sel_R_DATA_TEMPR105[24] ), 
        .C(sel_R_DATA_TEMPR106[24] ), .D(sel_R_DATA_TEMPR107[24] ), .Y(
        OR4_790_Y));
    OR4 OR4_1115 (.A(sel_R_DATA_TEMPR8[26] ), .B(sel_R_DATA_TEMPR9[26] ), .C(sel_R_DATA_TEMPR10[26] ), .D(sel_R_DATA_TEMPR11[26] ), .Y(OR4_1115_Y)
        );
    OR4 OR4_239 (.A(sel_R_DATA_TEMPR92[2] ), .B(sel_R_DATA_TEMPR93[2] ), .C(sel_R_DATA_TEMPR94[2] ), .D(sel_R_DATA_TEMPR95[2] ), .Y(OR4_239_Y));
    OR4 OR4_42 (.A(sel_R_DATA_TEMPR120[18] ), .B(sel_R_DATA_TEMPR121[18] ), 
        .C(sel_R_DATA_TEMPR122[18] ), .D(sel_R_DATA_TEMPR123[18] ), .Y(
        OR4_42_Y));
    OR4 OR4_529 (.A(sel_R_DATA_TEMPR108[31] ), .B(sel_R_DATA_TEMPR109[31] ), 
        .C(sel_R_DATA_TEMPR110[31] ), .D(sel_R_DATA_TEMPR111[31] ), .Y(
        OR4_529_Y));
    OR4 OR4_477 (.A(sel_R_DATA_TEMPR12[10] ), .B(sel_R_DATA_TEMPR13[10] ), 
        .C(sel_R_DATA_TEMPR14[10] ), .D(sel_R_DATA_TEMPR15[10] ), .Y(
        OR4_477_Y));
    OR4 OR4_1206 (.A(\DB_DETECT[104] ), .B(\DB_DETECT[105] ), .C(
        \DB_DETECT[106] ), .D(\DB_DETECT[107] ), .Y(OR4_1206_Y));
    OR4 OR4_1011 (.A(OR4_1362_Y), .B(OR4_229_Y), .C(OR4_444_Y), .D(
        OR4_279_Y), .Y(OR4_1011_Y));
    OR4 OR4_492 (.A(sel_R_DATA_TEMPR104[22] ), .B(sel_R_DATA_TEMPR105[22] ), 
        .C(sel_R_DATA_TEMPR106[22] ), .D(sel_R_DATA_TEMPR107[22] ), .Y(
        OR4_492_Y));
    AND4 \AND4SB_CORRECT[38]  (.A(sel_SB_CORRECT_NG[38] ), .B(
        \BLKY2_pipe[9] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[38] ));
    AND4 \AND4DB_DETECT[112]  (.A(sel_DB_DETECT_NG[112] ), .B(
        \BLKY2_pipe[28] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[112] ));
    AND4 \AND4DB_DETECT[4]  (.A(sel_DB_DETECT_NG[4] ), .B(
        \BLKY2_pipe[1] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[4] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%114%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R114C0 (.A_DOUT({
        nc248, nc249, nc250, nc251, nc252,int_R_DATA_TEMPR114[31] , 
       int_R_DATA_TEMPR114[30] ,int_R_DATA_TEMPR114[29] , 
       int_R_DATA_TEMPR114[28] ,int_R_DATA_TEMPR114[27] , 
       int_R_DATA_TEMPR114[26] ,int_R_DATA_TEMPR114[25] , 
       int_R_DATA_TEMPR114[24] ,int_R_DATA_TEMPR114[23] , 
       int_R_DATA_TEMPR114[22] ,int_R_DATA_TEMPR114[21] , 
       int_R_DATA_TEMPR114[20] ,int_R_DATA_TEMPR114[19] , 
       int_R_DATA_TEMPR114[18] ,int_R_DATA_TEMPR114[17] }), .B_DOUT({nc253, 
        nc254, nc255,int_R_DATA_TEMPR114[16] ,int_R_DATA_TEMPR114[15] , 
       int_R_DATA_TEMPR114[14] ,int_R_DATA_TEMPR114[13] , 
       int_R_DATA_TEMPR114[12] ,int_R_DATA_TEMPR114[11] , 
       int_R_DATA_TEMPR114[10] ,int_R_DATA_TEMPR114[9] , 
       int_R_DATA_TEMPR114[8] ,int_R_DATA_TEMPR114[7] , 
       int_R_DATA_TEMPR114[6] ,int_R_DATA_TEMPR114[5] , 
       int_R_DATA_TEMPR114[4] ,int_R_DATA_TEMPR114[3] , 
       int_R_DATA_TEMPR114[2] ,int_R_DATA_TEMPR114[1] , 
       int_R_DATA_TEMPR114[0] }), .DB_DETECT(int_DB_DETECT_NG[114] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[114] ), .ACCESS_BUSY(
        ACCESS_BUSY[114] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[28] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[28] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_520 (.A(sel_R_DATA_TEMPR44[12] ), .B(sel_R_DATA_TEMPR45[12] ), 
        .C(sel_R_DATA_TEMPR46[12] ), .D(sel_R_DATA_TEMPR47[12] ), .Y(
        OR4_520_Y));
    OR4 OR4_499 (.A(sel_R_DATA_TEMPR100[27] ), .B(sel_R_DATA_TEMPR101[27] ), 
        .C(sel_R_DATA_TEMPR102[27] ), .D(sel_R_DATA_TEMPR103[27] ), .Y(
        OR4_499_Y));
    OR4 OR4_88 (.A(sel_R_DATA_TEMPR0[20] ), .B(sel_R_DATA_TEMPR1[20] ), .C(sel_R_DATA_TEMPR2[20] ), .D(sel_R_DATA_TEMPR3[20] ), .Y(OR4_88_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[7]  (.A(CFG3_23_Y), .B(
        CFG3_12_Y), .Y(\BLKX2[7] ));
    OR4 OR4_1308 (.A(sel_R_DATA_TEMPR4[9] ), .B(sel_R_DATA_TEMPR5[9] ), .C(sel_R_DATA_TEMPR6[9] ), .D(sel_R_DATA_TEMPR7[9] ), .Y(OR4_1308_Y));
    OR4 OR4_205 (.A(sel_R_DATA_TEMPR24[10] ), .B(sel_R_DATA_TEMPR25[10] ), 
        .C(sel_R_DATA_TEMPR26[10] ), .D(sel_R_DATA_TEMPR27[10] ), .Y(
        OR4_205_Y));
    OR4 OR4_887 (.A(sel_R_DATA_TEMPR92[21] ), .B(sel_R_DATA_TEMPR93[21] ), 
        .C(sel_R_DATA_TEMPR94[21] ), .D(sel_R_DATA_TEMPR95[21] ), .Y(
        OR4_887_Y));
    AND4 \AND4DB_DETECT[85]  (.A(sel_DB_DETECT_NG[85] ), .B(
        \BLKY2_pipe[21] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[85] ));
    OR4 OR4_188 (.A(sel_R_DATA_TEMPR16[17] ), .B(sel_R_DATA_TEMPR17[17] ), 
        .C(sel_R_DATA_TEMPR18[17] ), .D(sel_R_DATA_TEMPR19[17] ), .Y(
        OR4_188_Y));
    OR4 OR4_984 (.A(sel_R_DATA_TEMPR96[8] ), .B(sel_R_DATA_TEMPR97[8] ), .C(sel_R_DATA_TEMPR98[8] ), .D(sel_R_DATA_TEMPR99[8] ), .Y(OR4_984_Y));
    OR4 OR4_810 (.A(\DB_DETECT[28] ), .B(\DB_DETECT[29] ), .C(
        \DB_DETECT[30] ), .D(\DB_DETECT[31] ), .Y(OR4_810_Y));
    OR4 OR4_196 (.A(sel_R_DATA_TEMPR116[20] ), .B(sel_R_DATA_TEMPR117[20] ), 
        .C(sel_R_DATA_TEMPR118[20] ), .D(sel_R_DATA_TEMPR119[20] ), .Y(
        OR4_196_Y));
    OR4 OR4_802 (.A(sel_R_DATA_TEMPR120[6] ), .B(sel_R_DATA_TEMPR121[6] ), 
        .C(sel_R_DATA_TEMPR122[6] ), .D(sel_R_DATA_TEMPR123[6] ), .Y(
        OR4_802_Y));
    OR4 OR4_112 (.A(sel_R_DATA_TEMPR32[16] ), .B(sel_R_DATA_TEMPR33[16] ), 
        .C(sel_R_DATA_TEMPR34[16] ), .D(sel_R_DATA_TEMPR35[16] ), .Y(
        OR4_112_Y));
    OR4 OR4_275 (.A(sel_R_DATA_TEMPR116[25] ), .B(sel_R_DATA_TEMPR117[25] ), 
        .C(sel_R_DATA_TEMPR118[25] ), .D(sel_R_DATA_TEMPR119[25] ), .Y(
        OR4_275_Y));
    OR4 OR4_1270 (.A(sel_R_DATA_TEMPR20[9] ), .B(sel_R_DATA_TEMPR21[9] ), .C(sel_R_DATA_TEMPR22[9] ), .D(sel_R_DATA_TEMPR23[9] ), .Y(OR4_1270_Y));
    OR4 OR4_1013 (.A(OR4_294_Y), .B(OR4_862_Y), .C(OR4_1343_Y), .D(
        OR4_813_Y), .Y(OR4_1013_Y));
    OR4 OR4_915 (.A(sel_R_DATA_TEMPR88[19] ), .B(sel_R_DATA_TEMPR89[19] ), 
        .C(sel_R_DATA_TEMPR90[19] ), .D(sel_R_DATA_TEMPR91[19] ), .Y(
        OR4_915_Y));
    OR4 OR4_839 (.A(sel_R_DATA_TEMPR100[26] ), .B(sel_R_DATA_TEMPR101[26] ), 
        .C(sel_R_DATA_TEMPR102[26] ), .D(sel_R_DATA_TEMPR103[26] ), .Y(
        OR4_839_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%107%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R107C0 (.A_DOUT({
        nc256, nc257, nc258, nc259, nc260,int_R_DATA_TEMPR107[31] , 
       int_R_DATA_TEMPR107[30] ,int_R_DATA_TEMPR107[29] , 
       int_R_DATA_TEMPR107[28] ,int_R_DATA_TEMPR107[27] , 
       int_R_DATA_TEMPR107[26] ,int_R_DATA_TEMPR107[25] , 
       int_R_DATA_TEMPR107[24] ,int_R_DATA_TEMPR107[23] , 
       int_R_DATA_TEMPR107[22] ,int_R_DATA_TEMPR107[21] , 
       int_R_DATA_TEMPR107[20] ,int_R_DATA_TEMPR107[19] , 
       int_R_DATA_TEMPR107[18] ,int_R_DATA_TEMPR107[17] }), .B_DOUT({nc261, 
        nc262, nc263,int_R_DATA_TEMPR107[16] ,int_R_DATA_TEMPR107[15] , 
       int_R_DATA_TEMPR107[14] ,int_R_DATA_TEMPR107[13] , 
       int_R_DATA_TEMPR107[12] ,int_R_DATA_TEMPR107[11] , 
       int_R_DATA_TEMPR107[10] ,int_R_DATA_TEMPR107[9] , 
       int_R_DATA_TEMPR107[8] ,int_R_DATA_TEMPR107[7] , 
       int_R_DATA_TEMPR107[6] ,int_R_DATA_TEMPR107[5] , 
       int_R_DATA_TEMPR107[4] ,int_R_DATA_TEMPR107[3] , 
       int_R_DATA_TEMPR107[2] ,int_R_DATA_TEMPR107[1] , 
       int_R_DATA_TEMPR107[0] }), .DB_DETECT(int_DB_DETECT_NG[107] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[107] ), .ACCESS_BUSY(
        ACCESS_BUSY[107] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[26] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[26] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4DB_DETECT[100]  (.A(sel_DB_DETECT_NG[100] ), .B(
        \BLKY2_pipe[25] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[100] ));
    OR4 OR4_872 (.A(sel_R_DATA_TEMPR100[6] ), .B(sel_R_DATA_TEMPR101[6] ), 
        .C(sel_R_DATA_TEMPR102[6] ), .D(sel_R_DATA_TEMPR103[6] ), .Y(
        OR4_872_Y));
    OR4 OR4_646 (.A(OR4_711_Y), .B(OR4_1216_Y), .C(OR4_492_Y), .D(
        OR4_696_Y), .Y(OR4_646_Y));
    AND4 \AND4SB_CORRECT[23]  (.A(sel_SB_CORRECT_NG[23] ), .B(
        \BLKY2_pipe[5] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[23] ));
    AND4 \AND4DB_DETECT[72]  (.A(sel_DB_DETECT_NG[72] ), .B(
        \BLKY2_pipe[18] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[72] ));
    OR4 OR4_1286 (.A(OR4_219_Y), .B(OR4_207_Y), .C(OR4_658_Y), .D(
        OR4_146_Y), .Y(OR4_1286_Y));
    OR4 OR4_257 (.A(sel_R_DATA_TEMPR36[20] ), .B(sel_R_DATA_TEMPR37[20] ), 
        .C(sel_R_DATA_TEMPR38[20] ), .D(sel_R_DATA_TEMPR39[20] ), .Y(
        OR4_257_Y));
    AND4 \AND4SB_CORRECT[19]  (.A(sel_SB_CORRECT_NG[19] ), .B(
        \BLKY2_pipe[4] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[19] ));
    OR4 OR4_1372 (.A(sel_R_DATA_TEMPR96[4] ), .B(sel_R_DATA_TEMPR97[4] ), .C(sel_R_DATA_TEMPR98[4] ), .D(sel_R_DATA_TEMPR99[4] ), .Y(OR4_1372_Y));
    OR4 OR4_398 (.A(sel_R_DATA_TEMPR64[16] ), .B(sel_R_DATA_TEMPR65[16] ), 
        .C(sel_R_DATA_TEMPR66[16] ), .D(sel_R_DATA_TEMPR67[16] ), .Y(
        OR4_398_Y));
    OR4 OR4_1009 (.A(sel_R_DATA_TEMPR124[6] ), .B(sel_R_DATA_TEMPR125[6] ), 
        .C(sel_R_DATA_TEMPR126[6] ), .D(sel_R_DATA_TEMPR127[6] ), .Y(
        OR4_1009_Y));
    OR4 OR4_157 (.A(sel_R_DATA_TEMPR100[10] ), .B(sel_R_DATA_TEMPR101[10] ), 
        .C(sel_R_DATA_TEMPR102[10] ), .D(sel_R_DATA_TEMPR103[10] ), .Y(
        OR4_157_Y));
    OR4 OR4_1335 (.A(\SB_CORRECT[44] ), .B(\SB_CORRECT[45] ), .C(
        \SB_CORRECT[46] ), .D(\SB_CORRECT[47] ), .Y(OR4_1335_Y));
    OR4 OR4_1272 (.A(OR4_374_Y), .B(OR4_829_Y), .C(OR4_1297_Y), .D(
        OR4_301_Y), .Y(OR4_1272_Y));
    OR4 OR4_561 (.A(OR4_717_Y), .B(OR4_938_Y), .C(OR4_1101_Y), .D(
        OR4_735_Y), .Y(OR4_561_Y));
    OR4 OR4_403 (.A(sel_R_DATA_TEMPR120[17] ), .B(sel_R_DATA_TEMPR121[17] ), 
        .C(sel_R_DATA_TEMPR122[17] ), .D(sel_R_DATA_TEMPR123[17] ), .Y(
        OR4_403_Y));
    OR4 OR4_1388 (.A(sel_R_DATA_TEMPR44[8] ), .B(sel_R_DATA_TEMPR45[8] ), .C(sel_R_DATA_TEMPR46[8] ), .D(sel_R_DATA_TEMPR47[8] ), .Y(OR4_1388_Y));
    OR4 OR4_1153 (.A(OR4_1226_Y), .B(OR2_7_Y), .C(sel_R_DATA_TEMPR86[1] ), 
        .D(sel_R_DATA_TEMPR87[1] ), .Y(OR4_1153_Y));
    OR4 OR4_601 (.A(sel_R_DATA_TEMPR124[31] ), .B(sel_R_DATA_TEMPR125[31] ), 
        .C(sel_R_DATA_TEMPR126[31] ), .D(sel_R_DATA_TEMPR127[31] ), .Y(
        OR4_601_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_7 (.A(W_EN), .B(W_ADDR[15]), .C(
        W_ADDR[14]), .Y(CFG3_7_Y));
    OR4 OR4_1164 (.A(sel_R_DATA_TEMPR64[15] ), .B(sel_R_DATA_TEMPR65[15] ), 
        .C(sel_R_DATA_TEMPR66[15] ), .D(sel_R_DATA_TEMPR67[15] ), .Y(
        OR4_1164_Y));
    OR4 OR4_208 (.A(sel_R_DATA_TEMPR8[10] ), .B(sel_R_DATA_TEMPR9[10] ), .C(sel_R_DATA_TEMPR10[10] ), .D(sel_R_DATA_TEMPR11[10] ), .Y(OR4_208_Y));
    OR4 OR4_219 (.A(OR4_924_Y), .B(OR4_698_Y), .C(OR4_471_Y), .D(
        OR4_1278_Y), .Y(OR4_219_Y));
    OR4 \OR4_R_DATA[19]  (.A(OR4_447_Y), .B(OR4_129_Y), .C(OR4_37_Y), 
        .D(OR4_1197_Y), .Y(R_DATA[19]));
    OR4 OR4_323 (.A(OR4_189_Y), .B(OR4_636_Y), .C(OR4_333_Y), .D(
        OR4_330_Y), .Y(OR4_323_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[19]  (.A(CFG3_19_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[19] ));
    OR4 OR4_720 (.A(OR4_79_Y), .B(OR4_1321_Y), .C(OR4_38_Y), .D(
        OR4_1339_Y), .Y(OR4_720_Y));
    OR4 OR4_473 (.A(sel_R_DATA_TEMPR4[6] ), .B(sel_R_DATA_TEMPR5[6] ), .C(sel_R_DATA_TEMPR6[6] ), .D(sel_R_DATA_TEMPR7[6] ), .Y(OR4_473_Y));
    AND4 \AND4DB_DETECT[110]  (.A(sel_DB_DETECT_NG[110] ), .B(
        \BLKY2_pipe[27] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[110] ));
    OR4 OR4_671 (.A(OR4_920_Y), .B(OR4_1140_Y), .C(OR4_1301_Y), .D(
        OR4_1296_Y), .Y(OR4_671_Y));
    OR4 OR4_737 (.A(sel_R_DATA_TEMPR8[9] ), .B(sel_R_DATA_TEMPR9[9] ), .C(sel_R_DATA_TEMPR10[9] ), .D(sel_R_DATA_TEMPR11[9] ), .Y(OR4_737_Y));
    OR4 OR4_422 (.A(sel_R_DATA_TEMPR0[5] ), .B(sel_R_DATA_TEMPR1[5] ), .C(sel_R_DATA_TEMPR2[5] ), .D(sel_R_DATA_TEMPR3[5] ), .Y(OR4_422_Y));
    OR4 OR4_278 (.A(sel_R_DATA_TEMPR44[22] ), .B(sel_R_DATA_TEMPR45[22] ), 
        .C(sel_R_DATA_TEMPR46[22] ), .D(sel_R_DATA_TEMPR47[22] ), .Y(
        OR4_278_Y));
    OR4 OR4_753 (.A(sel_R_DATA_TEMPR36[16] ), .B(sel_R_DATA_TEMPR37[16] ), 
        .C(sel_R_DATA_TEMPR38[16] ), .D(sel_R_DATA_TEMPR39[16] ), .Y(
        OR4_753_Y));
    OR4 OR4_734 (.A(sel_R_DATA_TEMPR116[27] ), .B(sel_R_DATA_TEMPR117[27] ), 
        .C(sel_R_DATA_TEMPR118[27] ), .D(sel_R_DATA_TEMPR119[27] ), .Y(
        OR4_734_Y));
    OR4 OR4_1274 (.A(sel_R_DATA_TEMPR36[12] ), .B(sel_R_DATA_TEMPR37[12] ), 
        .C(sel_R_DATA_TEMPR38[12] ), .D(sel_R_DATA_TEMPR39[12] ), .Y(
        OR4_1274_Y));
    AND4 \AND4SB_CORRECT[24]  (.A(sel_SB_CORRECT_NG[24] ), .B(
        \BLKY2_pipe[6] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[24] ));
    OR4 OR4_23 (.A(sel_R_DATA_TEMPR20[17] ), .B(sel_R_DATA_TEMPR21[17] ), .C(sel_R_DATA_TEMPR22[17] ), .D(sel_R_DATA_TEMPR23[17] ), .Y(OR4_23_Y));
    OR4 OR4_199 (.A(\DB_DETECT[32] ), .B(\DB_DETECT[33] ), .C(
        \DB_DETECT[34] ), .D(\DB_DETECT[35] ), .Y(OR4_199_Y));
    OR4 OR4_254 (.A(OR4_504_Y), .B(OR4_1379_Y), .C(OR4_194_Y), .D(
        OR4_675_Y), .Y(OR4_254_Y));
    AND4 \AND4DB_DETECT[29]  (.A(sel_DB_DETECT_NG[29] ), .B(
        \BLKY2_pipe[7] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[29] ));
    OR4 OR4_429 (.A(OR4_804_Y), .B(OR2_16_Y), .C(sel_R_DATA_TEMPR86[30] ), 
        .D(sel_R_DATA_TEMPR87[30] ), .Y(OR4_429_Y));
    OR4 OR4_1268 (.A(\SB_CORRECT[64] ), .B(\SB_CORRECT[65] ), .C(
        \SB_CORRECT[66] ), .D(\SB_CORRECT[67] ), .Y(OR4_1268_Y));
    OR4 OR4_262 (.A(sel_R_DATA_TEMPR44[18] ), .B(sel_R_DATA_TEMPR45[18] ), 
        .C(sel_R_DATA_TEMPR46[18] ), .D(sel_R_DATA_TEMPR47[18] ), .Y(
        OR4_262_Y));
    OR4 OR4_1377 (.A(sel_R_DATA_TEMPR12[17] ), .B(sel_R_DATA_TEMPR13[17] ), 
        .C(sel_R_DATA_TEMPR14[17] ), .D(sel_R_DATA_TEMPR15[17] ), .Y(
        OR4_1377_Y));
    AND4 \AND4SB_CORRECT[40]  (.A(sel_SB_CORRECT_NG[40] ), .B(
        \BLKY2_pipe[10] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[40] ));
    OR4 OR4_1249 (.A(OR4_1184_Y), .B(OR4_692_Y), .C(OR4_90_Y), .D(
        OR4_879_Y), .Y(OR4_1249_Y));
    OR4 OR4_1089 (.A(OR4_1307_Y), .B(OR4_575_Y), .C(OR4_968_Y), .D(
        OR4_1255_Y), .Y(OR4_1089_Y));
    OR4 OR4_831 (.A(OR4_643_Y), .B(OR4_1250_Y), .C(OR4_312_Y), .D(
        OR4_1191_Y), .Y(OR4_831_Y));
    AND4 \AND4SB_CORRECT[63]  (.A(sel_SB_CORRECT_NG[63] ), .B(
        \BLKY2_pipe[15] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[63] ));
    OR4 OR4_126 (.A(sel_R_DATA_TEMPR100[24] ), .B(sel_R_DATA_TEMPR101[24] ), 
        .C(sel_R_DATA_TEMPR102[24] ), .D(sel_R_DATA_TEMPR103[24] ), .Y(
        OR4_126_Y));
    OR4 OR4_819 (.A(sel_R_DATA_TEMPR76[16] ), .B(sel_R_DATA_TEMPR77[16] ), 
        .C(sel_R_DATA_TEMPR78[16] ), .D(sel_R_DATA_TEMPR79[16] ), .Y(
        OR4_819_Y));
    OR4 OR4_94 (.A(sel_R_DATA_TEMPR116[0] ), .B(sel_R_DATA_TEMPR117[0] ), .C(sel_R_DATA_TEMPR118[0] ), .D(sel_R_DATA_TEMPR119[0] ), .Y(OR4_94_Y));
    OR4 OR4_1018 (.A(OR4_1045_Y), .B(OR4_627_Y), .C(OR4_607_Y), .D(
        OR4_345_Y), .Y(OR4_1018_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%80%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R80C0 (.A_DOUT({
        nc264, nc265, nc266, nc267, nc268,int_R_DATA_TEMPR80[31] , 
       int_R_DATA_TEMPR80[30] ,int_R_DATA_TEMPR80[29] , 
       int_R_DATA_TEMPR80[28] ,int_R_DATA_TEMPR80[27] , 
       int_R_DATA_TEMPR80[26] ,int_R_DATA_TEMPR80[25] , 
       int_R_DATA_TEMPR80[24] ,int_R_DATA_TEMPR80[23] , 
       int_R_DATA_TEMPR80[22] ,int_R_DATA_TEMPR80[21] , 
       int_R_DATA_TEMPR80[20] ,int_R_DATA_TEMPR80[19] , 
       int_R_DATA_TEMPR80[18] ,int_R_DATA_TEMPR80[17] }), .B_DOUT({nc269, 
        nc270, nc271,int_R_DATA_TEMPR80[16] ,int_R_DATA_TEMPR80[15] , 
       int_R_DATA_TEMPR80[14] ,int_R_DATA_TEMPR80[13] , 
       int_R_DATA_TEMPR80[12] ,int_R_DATA_TEMPR80[11] , 
       int_R_DATA_TEMPR80[10] ,int_R_DATA_TEMPR80[9] ,int_R_DATA_TEMPR80[8] , 
       int_R_DATA_TEMPR80[7] ,int_R_DATA_TEMPR80[6] ,int_R_DATA_TEMPR80[5] , 
       int_R_DATA_TEMPR80[4] ,int_R_DATA_TEMPR80[3] ,int_R_DATA_TEMPR80[2] , 
       int_R_DATA_TEMPR80[1] ,int_R_DATA_TEMPR80[0] }), .DB_DETECT( int_DB_DETECT_NG[80] ), .SB_CORRECT(int_SB_CORRECT_NG[80] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[80] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[20] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_65 (.A(sel_R_DATA_TEMPR96[0] ), .B(sel_R_DATA_TEMPR97[0] ), .C(sel_R_DATA_TEMPR98[0] ), .D(sel_R_DATA_TEMPR99[0] ), .Y(OR4_65_Y));
    OR4 OR4_991 (.A(sel_R_DATA_TEMPR36[18] ), .B(sel_R_DATA_TEMPR37[18] ), 
        .C(sel_R_DATA_TEMPR38[18] ), .D(sel_R_DATA_TEMPR39[18] ), .Y(
        OR4_991_Y));
    AND4 \AND4SB_CORRECT[120]  (.A(sel_SB_CORRECT_NG[120] ), .B(
        \BLKY2_pipe[30] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[120] ));
    OR4 OR4_360 (.A(sel_R_DATA_TEMPR0[7] ), .B(sel_R_DATA_TEMPR1[7] ), .C(sel_R_DATA_TEMPR2[7] ), .D(sel_R_DATA_TEMPR3[7] ), .Y(OR4_360_Y));
    OR4 OR4_1325 (.A(OR4_342_Y), .B(OR4_508_Y), .C(OR4_484_Y), .D(
        OR4_1144_Y), .Y(OR4_1325_Y));
    OR4 OR4_355 (.A(\SB_CORRECT[24] ), .B(\SB_CORRECT[25] ), .C(
        \SB_CORRECT[26] ), .D(\SB_CORRECT[27] ), .Y(OR4_355_Y));
    OR4 OR4_1194 (.A(sel_R_DATA_TEMPR48[5] ), .B(sel_R_DATA_TEMPR49[5] ), .C(sel_R_DATA_TEMPR50[5] ), .D(sel_R_DATA_TEMPR51[5] ), .Y(OR4_1194_Y));
    OR4 OR4_328 (.A(OR4_215_Y), .B(OR4_690_Y), .C(OR4_1378_Y), .D(
        OR4_204_Y), .Y(OR4_328_Y));
    OR4 OR4_344 (.A(sel_R_DATA_TEMPR100[18] ), .B(sel_R_DATA_TEMPR101[18] ), 
        .C(sel_R_DATA_TEMPR102[18] ), .D(sel_R_DATA_TEMPR103[18] ), .Y(
        OR4_344_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%17%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R17C0 (.A_DOUT({
        nc272, nc273, nc274, nc275, nc276,int_R_DATA_TEMPR17[31] , 
       int_R_DATA_TEMPR17[30] ,int_R_DATA_TEMPR17[29] , 
       int_R_DATA_TEMPR17[28] ,int_R_DATA_TEMPR17[27] , 
       int_R_DATA_TEMPR17[26] ,int_R_DATA_TEMPR17[25] , 
       int_R_DATA_TEMPR17[24] ,int_R_DATA_TEMPR17[23] , 
       int_R_DATA_TEMPR17[22] ,int_R_DATA_TEMPR17[21] , 
       int_R_DATA_TEMPR17[20] ,int_R_DATA_TEMPR17[19] , 
       int_R_DATA_TEMPR17[18] ,int_R_DATA_TEMPR17[17] }), .B_DOUT({nc277, 
        nc278, nc279,int_R_DATA_TEMPR17[16] ,int_R_DATA_TEMPR17[15] , 
       int_R_DATA_TEMPR17[14] ,int_R_DATA_TEMPR17[13] , 
       int_R_DATA_TEMPR17[12] ,int_R_DATA_TEMPR17[11] , 
       int_R_DATA_TEMPR17[10] ,int_R_DATA_TEMPR17[9] ,int_R_DATA_TEMPR17[8] , 
       int_R_DATA_TEMPR17[7] ,int_R_DATA_TEMPR17[6] ,int_R_DATA_TEMPR17[5] , 
       int_R_DATA_TEMPR17[4] ,int_R_DATA_TEMPR17[3] ,int_R_DATA_TEMPR17[2] , 
       int_R_DATA_TEMPR17[1] ,int_R_DATA_TEMPR17[0] }), .DB_DETECT( int_DB_DETECT_NG[17] ), .SB_CORRECT(int_SB_CORRECT_NG[17] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[17] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%118%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R118C0 (.A_DOUT({
        nc280, nc281, nc282, nc283, nc284,int_R_DATA_TEMPR118[31] , 
       int_R_DATA_TEMPR118[30] ,int_R_DATA_TEMPR118[29] , 
       int_R_DATA_TEMPR118[28] ,int_R_DATA_TEMPR118[27] , 
       int_R_DATA_TEMPR118[26] ,int_R_DATA_TEMPR118[25] , 
       int_R_DATA_TEMPR118[24] ,int_R_DATA_TEMPR118[23] , 
       int_R_DATA_TEMPR118[22] ,int_R_DATA_TEMPR118[21] , 
       int_R_DATA_TEMPR118[20] ,int_R_DATA_TEMPR118[19] , 
       int_R_DATA_TEMPR118[18] ,int_R_DATA_TEMPR118[17] }), .B_DOUT({nc285, 
        nc286, nc287,int_R_DATA_TEMPR118[16] ,int_R_DATA_TEMPR118[15] , 
       int_R_DATA_TEMPR118[14] ,int_R_DATA_TEMPR118[13] , 
       int_R_DATA_TEMPR118[12] ,int_R_DATA_TEMPR118[11] , 
       int_R_DATA_TEMPR118[10] ,int_R_DATA_TEMPR118[9] , 
       int_R_DATA_TEMPR118[8] ,int_R_DATA_TEMPR118[7] , 
       int_R_DATA_TEMPR118[6] ,int_R_DATA_TEMPR118[5] , 
       int_R_DATA_TEMPR118[4] ,int_R_DATA_TEMPR118[3] , 
       int_R_DATA_TEMPR118[2] ,int_R_DATA_TEMPR118[1] , 
       int_R_DATA_TEMPR118[0] }), .DB_DETECT(int_DB_DETECT_NG[118] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[118] ), .ACCESS_BUSY(
        ACCESS_BUSY[118] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[29] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[29] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_863 (.A(sel_R_DATA_TEMPR68[23] ), .B(sel_R_DATA_TEMPR69[23] ), 
        .C(sel_R_DATA_TEMPR70[23] ), .D(sel_R_DATA_TEMPR71[23] ), .Y(
        OR4_863_Y));
    OR4 OR4_185 (.A(sel_R_DATA_TEMPR20[23] ), .B(sel_R_DATA_TEMPR21[23] ), 
        .C(sel_R_DATA_TEMPR22[23] ), .D(sel_R_DATA_TEMPR23[23] ), .Y(
        OR4_185_Y));
    AND4 \AND4SB_CORRECT[64]  (.A(sel_SB_CORRECT_NG[64] ), .B(
        \BLKY2_pipe[16] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[64] ));
    OR4 OR4_141 (.A(sel_R_DATA_TEMPR112[11] ), .B(sel_R_DATA_TEMPR113[11] ), 
        .C(sel_R_DATA_TEMPR114[11] ), .D(sel_R_DATA_TEMPR115[11] ), .Y(
        OR4_141_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[16]  (.A(CFG3_16_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[16] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%76%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R76C0 (.A_DOUT({
        nc288, nc289, nc290, nc291, nc292,int_R_DATA_TEMPR76[31] , 
       int_R_DATA_TEMPR76[30] ,int_R_DATA_TEMPR76[29] , 
       int_R_DATA_TEMPR76[28] ,int_R_DATA_TEMPR76[27] , 
       int_R_DATA_TEMPR76[26] ,int_R_DATA_TEMPR76[25] , 
       int_R_DATA_TEMPR76[24] ,int_R_DATA_TEMPR76[23] , 
       int_R_DATA_TEMPR76[22] ,int_R_DATA_TEMPR76[21] , 
       int_R_DATA_TEMPR76[20] ,int_R_DATA_TEMPR76[19] , 
       int_R_DATA_TEMPR76[18] ,int_R_DATA_TEMPR76[17] }), .B_DOUT({nc293, 
        nc294, nc295,int_R_DATA_TEMPR76[16] ,int_R_DATA_TEMPR76[15] , 
       int_R_DATA_TEMPR76[14] ,int_R_DATA_TEMPR76[13] , 
       int_R_DATA_TEMPR76[12] ,int_R_DATA_TEMPR76[11] , 
       int_R_DATA_TEMPR76[10] ,int_R_DATA_TEMPR76[9] ,int_R_DATA_TEMPR76[8] , 
       int_R_DATA_TEMPR76[7] ,int_R_DATA_TEMPR76[6] ,int_R_DATA_TEMPR76[5] , 
       int_R_DATA_TEMPR76[4] ,int_R_DATA_TEMPR76[3] ,int_R_DATA_TEMPR76[2] , 
       int_R_DATA_TEMPR76[1] ,int_R_DATA_TEMPR76[0] }), .DB_DETECT( int_DB_DETECT_NG[76] ), .SB_CORRECT(int_SB_CORRECT_NG[76] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[76] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[19] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[19] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_717 (.A(sel_R_DATA_TEMPR64[3] ), .B(sel_R_DATA_TEMPR65[3] ), .C(sel_R_DATA_TEMPR66[3] ), .D(sel_R_DATA_TEMPR67[3] ), .Y(OR4_717_Y));
    OR4 OR4_36 (.A(sel_R_DATA_TEMPR96[1] ), .B(sel_R_DATA_TEMPR97[1] ), .C(sel_R_DATA_TEMPR98[1] ), .D(sel_R_DATA_TEMPR99[1] ), .Y(OR4_36_Y));
    OR4 OR4_487 (.A(sel_R_DATA_TEMPR28[15] ), .B(sel_R_DATA_TEMPR29[15] ), 
        .C(sel_R_DATA_TEMPR30[15] ), .D(sel_R_DATA_TEMPR31[15] ), .Y(
        OR4_487_Y));
    OR4 OR4_714 (.A(OR4_909_Y), .B(OR4_1128_Y), .C(OR4_1294_Y), .D(
        OR4_1099_Y), .Y(OR4_714_Y));
    OR4 OR4_501 (.A(sel_R_DATA_TEMPR108[4] ), .B(sel_R_DATA_TEMPR109[4] ), 
        .C(sel_R_DATA_TEMPR110[4] ), .D(sel_R_DATA_TEMPR111[4] ), .Y(
        OR4_501_Y));
    AND4 \AND4DB_DETECT[126]  (.A(sel_DB_DETECT_NG[126] ), .B(
        \BLKY2_pipe[31] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[126] ));
    CFG3 #( .INIT(8'h80) )  CFG3_23 (.A(W_ADDR[13]), .B(W_ADDR[12]), 
        .C(W_ADDR[11]), .Y(CFG3_23_Y));
    OR4 OR4_21 (.A(sel_R_DATA_TEMPR88[21] ), .B(sel_R_DATA_TEMPR89[21] ), .C(sel_R_DATA_TEMPR90[21] ), .D(sel_R_DATA_TEMPR91[21] ), .Y(OR4_21_Y));
    OR4 OR4_1298 (.A(sel_R_DATA_TEMPR116[23] ), .B(sel_R_DATA_TEMPR117[23] ), 
        .C(sel_R_DATA_TEMPR118[23] ), .D(sel_R_DATA_TEMPR119[23] ), .Y(
        OR4_1298_Y));
    OR4 OR4_1165 (.A(sel_R_DATA_TEMPR12[27] ), .B(sel_R_DATA_TEMPR13[27] ), 
        .C(sel_R_DATA_TEMPR14[27] ), .D(sel_R_DATA_TEMPR15[27] ), .Y(
        OR4_1165_Y));
    OR4 OR4_1107 (.A(sel_R_DATA_TEMPR48[9] ), .B(sel_R_DATA_TEMPR49[9] ), .C(sel_R_DATA_TEMPR50[9] ), .D(sel_R_DATA_TEMPR51[9] ), .Y(OR4_1107_Y));
    OR4 OR4_937 (.A(OR4_394_Y), .B(OR2_22_Y), .C(\SB_CORRECT[86] ), 
        .D(\SB_CORRECT[87] ), .Y(OR4_937_Y));
    OR4 OR4_1032 (.A(sel_R_DATA_TEMPR8[21] ), .B(sel_R_DATA_TEMPR9[21] ), .C(sel_R_DATA_TEMPR10[21] ), .D(sel_R_DATA_TEMPR11[21] ), .Y(OR4_1032_Y)
        );
    OR4 OR4_129 (.A(OR4_731_Y), .B(OR4_936_Y), .C(OR4_915_Y), .D(
        OR4_190_Y), .Y(OR4_129_Y));
    OR4 OR4_571 (.A(sel_R_DATA_TEMPR36[25] ), .B(sel_R_DATA_TEMPR37[25] ), 
        .C(sel_R_DATA_TEMPR38[25] ), .D(sel_R_DATA_TEMPR39[25] ), .Y(
        OR4_571_Y));
    OR4 OR4_1061 (.A(OR4_306_Y), .B(OR4_516_Y), .C(OR4_666_Y), .D(
        OR4_475_Y), .Y(OR4_1061_Y));
    OR4 OR4_811 (.A(sel_R_DATA_TEMPR120[3] ), .B(sel_R_DATA_TEMPR121[3] ), 
        .C(sel_R_DATA_TEMPR122[3] ), .D(sel_R_DATA_TEMPR123[3] ), .Y(
        OR4_811_Y));
    AND4 \AND4DB_DETECT[101]  (.A(sel_DB_DETECT_NG[101] ), .B(
        \BLKY2_pipe[25] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[101] ));
    OR4 OR4_1256 (.A(sel_R_DATA_TEMPR120[10] ), .B(sel_R_DATA_TEMPR121[10] ), 
        .C(sel_R_DATA_TEMPR122[10] ), .D(sel_R_DATA_TEMPR123[10] ), .Y(
        OR4_1256_Y));
    OR4 OR4_752 (.A(OR4_898_Y), .B(OR4_427_Y), .C(OR4_906_Y), .D(
        OR4_379_Y), .Y(OR4_752_Y));
    OR4 OR4_441 (.A(OR4_921_Y), .B(OR4_1308_Y), .C(OR4_737_Y), .D(
        OR4_995_Y), .Y(OR4_441_Y));
    OR4 OR4_795 (.A(sel_R_DATA_TEMPR16[21] ), .B(sel_R_DATA_TEMPR17[21] ), 
        .C(sel_R_DATA_TEMPR18[21] ), .D(sel_R_DATA_TEMPR19[21] ), .Y(
        OR4_795_Y));
    OR4 OR4_697 (.A(sel_R_DATA_TEMPR72[28] ), .B(sel_R_DATA_TEMPR73[28] ), 
        .C(sel_R_DATA_TEMPR74[28] ), .D(sel_R_DATA_TEMPR75[28] ), .Y(
        OR4_697_Y));
    AND4 \AND4SB_CORRECT[8]  (.A(sel_SB_CORRECT_NG[8] ), .B(
        \BLKY2_pipe[2] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[8] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%48%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R48C0 (.A_DOUT({
        nc296, nc297, nc298, nc299, nc300,int_R_DATA_TEMPR48[31] , 
       int_R_DATA_TEMPR48[30] ,int_R_DATA_TEMPR48[29] , 
       int_R_DATA_TEMPR48[28] ,int_R_DATA_TEMPR48[27] , 
       int_R_DATA_TEMPR48[26] ,int_R_DATA_TEMPR48[25] , 
       int_R_DATA_TEMPR48[24] ,int_R_DATA_TEMPR48[23] , 
       int_R_DATA_TEMPR48[22] ,int_R_DATA_TEMPR48[21] , 
       int_R_DATA_TEMPR48[20] ,int_R_DATA_TEMPR48[19] , 
       int_R_DATA_TEMPR48[18] ,int_R_DATA_TEMPR48[17] }), .B_DOUT({nc301, 
        nc302, nc303,int_R_DATA_TEMPR48[16] ,int_R_DATA_TEMPR48[15] , 
       int_R_DATA_TEMPR48[14] ,int_R_DATA_TEMPR48[13] , 
       int_R_DATA_TEMPR48[12] ,int_R_DATA_TEMPR48[11] , 
       int_R_DATA_TEMPR48[10] ,int_R_DATA_TEMPR48[9] ,int_R_DATA_TEMPR48[8] , 
       int_R_DATA_TEMPR48[7] ,int_R_DATA_TEMPR48[6] ,int_R_DATA_TEMPR48[5] , 
       int_R_DATA_TEMPR48[4] ,int_R_DATA_TEMPR48[3] ,int_R_DATA_TEMPR48[2] , 
       int_R_DATA_TEMPR48[1] ,int_R_DATA_TEMPR48[0] }), .DB_DETECT( int_DB_DETECT_NG[48] ), .SB_CORRECT(int_SB_CORRECT_NG[48] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[48] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[12] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[12] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_448 (.A(sel_R_DATA_TEMPR96[17] ), .B(sel_R_DATA_TEMPR97[17] ), 
        .C(sel_R_DATA_TEMPR98[17] ), .D(sel_R_DATA_TEMPR99[17] ), .Y(
        OR4_448_Y));
    OR4 OR4_796 (.A(sel_R_DATA_TEMPR88[6] ), .B(sel_R_DATA_TEMPR89[6] ), .C(sel_R_DATA_TEMPR90[6] ), .D(sel_R_DATA_TEMPR91[6] ), .Y(OR4_796_Y));
    OR4 OR4_285 (.A(sel_R_DATA_TEMPR108[30] ), .B(sel_R_DATA_TEMPR109[30] ), 
        .C(sel_R_DATA_TEMPR110[30] ), .D(sel_R_DATA_TEMPR111[30] ), .Y(
        OR4_285_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%45%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R45C0 (.A_DOUT({
        nc304, nc305, nc306, nc307, nc308,int_R_DATA_TEMPR45[31] , 
       int_R_DATA_TEMPR45[30] ,int_R_DATA_TEMPR45[29] , 
       int_R_DATA_TEMPR45[28] ,int_R_DATA_TEMPR45[27] , 
       int_R_DATA_TEMPR45[26] ,int_R_DATA_TEMPR45[25] , 
       int_R_DATA_TEMPR45[24] ,int_R_DATA_TEMPR45[23] , 
       int_R_DATA_TEMPR45[22] ,int_R_DATA_TEMPR45[21] , 
       int_R_DATA_TEMPR45[20] ,int_R_DATA_TEMPR45[19] , 
       int_R_DATA_TEMPR45[18] ,int_R_DATA_TEMPR45[17] }), .B_DOUT({nc309, 
        nc310, nc311,int_R_DATA_TEMPR45[16] ,int_R_DATA_TEMPR45[15] , 
       int_R_DATA_TEMPR45[14] ,int_R_DATA_TEMPR45[13] , 
       int_R_DATA_TEMPR45[12] ,int_R_DATA_TEMPR45[11] , 
       int_R_DATA_TEMPR45[10] ,int_R_DATA_TEMPR45[9] ,int_R_DATA_TEMPR45[8] , 
       int_R_DATA_TEMPR45[7] ,int_R_DATA_TEMPR45[6] ,int_R_DATA_TEMPR45[5] , 
       int_R_DATA_TEMPR45[4] ,int_R_DATA_TEMPR45[3] ,int_R_DATA_TEMPR45[2] , 
       int_R_DATA_TEMPR45[1] ,int_R_DATA_TEMPR45[0] }), .DB_DETECT( int_DB_DETECT_NG[45] ), .SB_CORRECT(int_SB_CORRECT_NG[45] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[45] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[11] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1358 (.A(sel_R_DATA_TEMPR60[26] ), .B(sel_R_DATA_TEMPR61[26] ), 
        .C(sel_R_DATA_TEMPR62[26] ), .D(sel_R_DATA_TEMPR63[26] ), .Y(
        OR4_1358_Y));
    OR4 OR4_956 (.A(sel_R_DATA_TEMPR28[12] ), .B(sel_R_DATA_TEMPR29[12] ), 
        .C(sel_R_DATA_TEMPR30[12] ), .D(sel_R_DATA_TEMPR31[12] ), .Y(
        OR4_956_Y));
    OR4 OR4_882 (.A(sel_R_DATA_TEMPR108[19] ), .B(sel_R_DATA_TEMPR109[19] ), 
        .C(sel_R_DATA_TEMPR110[19] ), .D(sel_R_DATA_TEMPR111[19] ), .Y(
        OR4_882_Y));
    OR4 OR4_202 (.A(OR4_1368_Y), .B(OR4_689_Y), .C(OR4_1386_Y), .D(
        OR4_212_Y), .Y(OR4_202_Y));
    OR4 OR4_655 (.A(sel_R_DATA_TEMPR116[3] ), .B(sel_R_DATA_TEMPR117[3] ), 
        .C(sel_R_DATA_TEMPR118[3] ), .D(sel_R_DATA_TEMPR119[3] ), .Y(
        OR4_655_Y));
    OR4 OR4_921 (.A(sel_R_DATA_TEMPR0[9] ), .B(sel_R_DATA_TEMPR1[9] ), .C(sel_R_DATA_TEMPR2[9] ), .D(sel_R_DATA_TEMPR3[9] ), .Y(OR4_921_Y));
    AND4 \AND4DB_DETECT[53]  (.A(sel_DB_DETECT_NG[53] ), .B(
        \BLKY2_pipe[13] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[53] ));
    OR4 OR4_1063 (.A(sel_R_DATA_TEMPR36[24] ), .B(sel_R_DATA_TEMPR37[24] ), 
        .C(sel_R_DATA_TEMPR38[24] ), .D(sel_R_DATA_TEMPR39[24] ), .Y(
        OR4_1063_Y));
    CFG3 #( .INIT(8'h1) )  CFG3_13 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_13_Y));
    AND4 \AND4SB_CORRECT[1]  (.A(sel_SB_CORRECT_NG[1] ), .B(
        \BLKY2_pipe[0] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[1] ));
    AND4 \AND4SB_CORRECT[85]  (.A(sel_SB_CORRECT_NG[85] ), .B(
        \BLKY2_pipe[21] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[85] ));
    AND4 \AND4SB_CORRECT[86]  (.A(sel_SB_CORRECT_NG[86] ), .B(
        \BLKY2_pipe[21] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[86] ));
    OR4 OR4_272 (.A(OR4_105_Y), .B(OR4_1085_Y), .C(OR4_156_Y), .D(
        OR4_540_Y), .Y(OR4_272_Y));
    AND4 \AND4DB_DETECT[44]  (.A(sel_DB_DETECT_NG[44] ), .B(
        \BLKY2_pipe[11] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[44] ));
    OR4 OR4_1187 (.A(sel_R_DATA_TEMPR32[30] ), .B(sel_R_DATA_TEMPR33[30] ), 
        .C(sel_R_DATA_TEMPR34[30] ), .D(sel_R_DATA_TEMPR35[30] ), .Y(
        OR4_1187_Y));
    OR4 OR4_1017 (.A(sel_R_DATA_TEMPR108[24] ), .B(sel_R_DATA_TEMPR109[24] ), 
        .C(sel_R_DATA_TEMPR110[24] ), .D(sel_R_DATA_TEMPR111[24] ), .Y(
        OR4_1017_Y));
    AND4 \AND4DB_DETECT[111]  (.A(sel_DB_DETECT_NG[111] ), .B(
        \BLKY2_pipe[27] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[111] ));
    OR4 OR4_1376 (.A(sel_R_DATA_TEMPR40[7] ), .B(sel_R_DATA_TEMPR41[7] ), .C(sel_R_DATA_TEMPR42[7] ), .D(sel_R_DATA_TEMPR43[7] ), .Y(OR4_1376_Y));
    OR4 OR4_565 (.A(sel_R_DATA_TEMPR64[13] ), .B(sel_R_DATA_TEMPR65[13] ), 
        .C(sel_R_DATA_TEMPR66[13] ), .D(sel_R_DATA_TEMPR67[13] ), .Y(
        OR4_565_Y));
    OR4 OR4_44 (.A(OR4_424_Y), .B(OR4_196_Y), .C(OR4_1349_Y), .D(
        OR4_1001_Y), .Y(OR4_44_Y));
    OR4 OR4_549 (.A(sel_R_DATA_TEMPR16[11] ), .B(sel_R_DATA_TEMPR17[11] ), 
        .C(sel_R_DATA_TEMPR18[11] ), .D(sel_R_DATA_TEMPR19[11] ), .Y(
        OR4_549_Y));
    AND4 \AND4DB_DETECT[103]  (.A(sel_DB_DETECT_NG[103] ), .B(
        \BLKY2_pipe[25] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[103] ));
    OR4 OR4_435 (.A(OR4_982_Y), .B(OR4_1265_Y), .C(OR4_82_Y), .D(
        OR4_1300_Y), .Y(OR4_435_Y));
    OR4 OR4_300 (.A(sel_R_DATA_TEMPR20[8] ), .B(sel_R_DATA_TEMPR21[8] ), .C(sel_R_DATA_TEMPR22[8] ), .D(sel_R_DATA_TEMPR23[8] ), .Y(OR4_300_Y));
    OR4 OR4_540 (.A(sel_R_DATA_TEMPR92[4] ), .B(sel_R_DATA_TEMPR93[4] ), .C(sel_R_DATA_TEMPR94[4] ), .D(sel_R_DATA_TEMPR95[4] ), .Y(OR4_540_Y));
    OR4 OR4_483 (.A(sel_R_DATA_TEMPR48[22] ), .B(sel_R_DATA_TEMPR49[22] ), 
        .C(sel_R_DATA_TEMPR50[22] ), .D(sel_R_DATA_TEMPR51[22] ), .Y(
        OR4_483_Y));
    OR4 OR4_1243 (.A(sel_R_DATA_TEMPR20[29] ), .B(sel_R_DATA_TEMPR21[29] ), 
        .C(sel_R_DATA_TEMPR22[29] ), .D(sel_R_DATA_TEMPR23[29] ), .Y(
        OR4_1243_Y));
    OR4 OR4_1059 (.A(sel_R_DATA_TEMPR44[17] ), .B(sel_R_DATA_TEMPR45[17] ), 
        .C(sel_R_DATA_TEMPR46[17] ), .D(sel_R_DATA_TEMPR47[17] ), .Y(
        OR4_1059_Y));
    OR4 OR4_681 (.A(sel_R_DATA_TEMPR32[23] ), .B(sel_R_DATA_TEMPR33[23] ), 
        .C(sel_R_DATA_TEMPR34[23] ), .D(sel_R_DATA_TEMPR35[23] ), .Y(
        OR4_681_Y));
    OR4 OR4_663 (.A(\SB_CORRECT[76] ), .B(\SB_CORRECT[77] ), .C(
        \SB_CORRECT[78] ), .D(\SB_CORRECT[79] ), .Y(OR4_663_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[22]  (.A(CFG3_1_Y), .B(CFG3_9_Y)
        , .Y(\BLKY2[22] ));
    OR4 OR4_1195 (.A(sel_R_DATA_TEMPR48[7] ), .B(sel_R_DATA_TEMPR49[7] ), .C(sel_R_DATA_TEMPR50[7] ), .D(sel_R_DATA_TEMPR51[7] ), .Y(OR4_1195_Y));
    OR4 OR4_370 (.A(sel_R_DATA_TEMPR52[11] ), .B(sel_R_DATA_TEMPR53[11] ), 
        .C(sel_R_DATA_TEMPR54[11] ), .D(sel_R_DATA_TEMPR55[11] ), .Y(
        OR4_370_Y));
    OR4 OR4_288 (.A(OR4_826_Y), .B(OR4_1103_Y), .C(OR4_1304_Y), .D(
        OR4_1141_Y), .Y(OR4_288_Y));
    OR4 OR4_917 (.A(\SB_CORRECT[40] ), .B(\SB_CORRECT[41] ), .C(
        \SB_CORRECT[42] ), .D(\SB_CORRECT[43] ), .Y(OR4_917_Y));
    CFG3 #( .INIT(8'h4) )  CFG3_0 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_0_Y));
    OR4 OR4_1022 (.A(sel_R_DATA_TEMPR20[21] ), .B(sel_R_DATA_TEMPR21[21] ), 
        .C(sel_R_DATA_TEMPR22[21] ), .D(sel_R_DATA_TEMPR23[21] ), .Y(
        OR4_1022_Y));
    AND4 \AND4SB_CORRECT[37]  (.A(sel_SB_CORRECT_NG[37] ), .B(
        \BLKY2_pipe[9] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[37] ));
    OR4 OR4_1091 (.A(sel_R_DATA_TEMPR40[3] ), .B(sel_R_DATA_TEMPR41[3] ), .C(sel_R_DATA_TEMPR42[3] ), .D(sel_R_DATA_TEMPR43[3] ), .Y(OR4_1091_Y));
    OR4 OR4_803 (.A(sel_R_DATA_TEMPR88[3] ), .B(sel_R_DATA_TEMPR89[3] ), .C(sel_R_DATA_TEMPR90[3] ), .D(sel_R_DATA_TEMPR91[3] ), .Y(OR4_803_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%21%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R21C0 (.A_DOUT({
        nc312, nc313, nc314, nc315, nc316,int_R_DATA_TEMPR21[31] , 
       int_R_DATA_TEMPR21[30] ,int_R_DATA_TEMPR21[29] , 
       int_R_DATA_TEMPR21[28] ,int_R_DATA_TEMPR21[27] , 
       int_R_DATA_TEMPR21[26] ,int_R_DATA_TEMPR21[25] , 
       int_R_DATA_TEMPR21[24] ,int_R_DATA_TEMPR21[23] , 
       int_R_DATA_TEMPR21[22] ,int_R_DATA_TEMPR21[21] , 
       int_R_DATA_TEMPR21[20] ,int_R_DATA_TEMPR21[19] , 
       int_R_DATA_TEMPR21[18] ,int_R_DATA_TEMPR21[17] }), .B_DOUT({nc317, 
        nc318, nc319,int_R_DATA_TEMPR21[16] ,int_R_DATA_TEMPR21[15] , 
       int_R_DATA_TEMPR21[14] ,int_R_DATA_TEMPR21[13] , 
       int_R_DATA_TEMPR21[12] ,int_R_DATA_TEMPR21[11] , 
       int_R_DATA_TEMPR21[10] ,int_R_DATA_TEMPR21[9] ,int_R_DATA_TEMPR21[8] , 
       int_R_DATA_TEMPR21[7] ,int_R_DATA_TEMPR21[6] ,int_R_DATA_TEMPR21[5] , 
       int_R_DATA_TEMPR21[4] ,int_R_DATA_TEMPR21[3] ,int_R_DATA_TEMPR21[2] , 
       int_R_DATA_TEMPR21[1] ,int_R_DATA_TEMPR21[0] }), .DB_DETECT( int_DB_DETECT_NG[21] ), .SB_CORRECT(int_SB_CORRECT_NG[21] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[21] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[5] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1200 (.A(sel_R_DATA_TEMPR36[10] ), .B(sel_R_DATA_TEMPR37[10] ), 
        .C(sel_R_DATA_TEMPR38[10] ), .D(sel_R_DATA_TEMPR39[10] ), .Y(
        OR4_1200_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[8]  (.A(CFG3_16_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[8] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[12]  (.A(CFG3_6_Y), .B(CFG3_4_Y)
        , .Y(\BLKX2[12] ));
    AND4 \AND4SB_CORRECT[18]  (.A(sel_SB_CORRECT_NG[18] ), .B(
        \BLKY2_pipe[4] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[18] ));
    OR4 OR4_30 (.A(sel_R_DATA_TEMPR0[26] ), .B(sel_R_DATA_TEMPR1[26] ), .C(sel_R_DATA_TEMPR2[26] ), .D(sel_R_DATA_TEMPR3[26] ), .Y(OR4_30_Y));
    OR4 OR4_650 (.A(OR4_1002_Y), .B(OR4_1058_Y), .C(OR4_775_Y), .D(
        OR4_842_Y), .Y(OR4_650_Y));
    AND4 \AND4DB_DETECT[113]  (.A(sel_DB_DETECT_NG[113] ), .B(
        \BLKY2_pipe[28] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[113] ));
    OR4 OR4_873 (.A(OR4_1136_Y), .B(OR4_562_Y), .C(OR4_847_Y), .D(
        OR4_162_Y), .Y(OR4_873_Y));
    OR4 OR4_725 (.A(sel_R_DATA_TEMPR20[1] ), .B(sel_R_DATA_TEMPR21[1] ), .C(sel_R_DATA_TEMPR22[1] ), .D(sel_R_DATA_TEMPR23[1] ), .Y(OR4_725_Y));
    OR4 OR4_627 (.A(sel_R_DATA_TEMPR36[31] ), .B(sel_R_DATA_TEMPR37[31] ), 
        .C(sel_R_DATA_TEMPR38[31] ), .D(sel_R_DATA_TEMPR39[31] ), .Y(
        OR4_627_Y));
    OR4 OR4_297 (.A(OR4_945_Y), .B(OR4_300_Y), .C(OR4_959_Y), .D(
        OR4_1196_Y), .Y(OR4_297_Y));
    OR4 OR4_726 (.A(sel_R_DATA_TEMPR48[25] ), .B(sel_R_DATA_TEMPR49[25] ), 
        .C(sel_R_DATA_TEMPR50[25] ), .D(sel_R_DATA_TEMPR51[25] ), .Y(
        OR4_726_Y));
    OR4 OR4_37 (.A(OR4_574_Y), .B(OR4_840_Y), .C(OR4_1051_Y), .D(
        OR4_882_Y), .Y(OR4_37_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%69%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R69C0 (.A_DOUT({
        nc320, nc321, nc322, nc323, nc324,int_R_DATA_TEMPR69[31] , 
       int_R_DATA_TEMPR69[30] ,int_R_DATA_TEMPR69[29] , 
       int_R_DATA_TEMPR69[28] ,int_R_DATA_TEMPR69[27] , 
       int_R_DATA_TEMPR69[26] ,int_R_DATA_TEMPR69[25] , 
       int_R_DATA_TEMPR69[24] ,int_R_DATA_TEMPR69[23] , 
       int_R_DATA_TEMPR69[22] ,int_R_DATA_TEMPR69[21] , 
       int_R_DATA_TEMPR69[20] ,int_R_DATA_TEMPR69[19] , 
       int_R_DATA_TEMPR69[18] ,int_R_DATA_TEMPR69[17] }), .B_DOUT({nc325, 
        nc326, nc327,int_R_DATA_TEMPR69[16] ,int_R_DATA_TEMPR69[15] , 
       int_R_DATA_TEMPR69[14] ,int_R_DATA_TEMPR69[13] , 
       int_R_DATA_TEMPR69[12] ,int_R_DATA_TEMPR69[11] , 
       int_R_DATA_TEMPR69[10] ,int_R_DATA_TEMPR69[9] ,int_R_DATA_TEMPR69[8] , 
       int_R_DATA_TEMPR69[7] ,int_R_DATA_TEMPR69[6] ,int_R_DATA_TEMPR69[5] , 
       int_R_DATA_TEMPR69[4] ,int_R_DATA_TEMPR69[3] ,int_R_DATA_TEMPR69[2] , 
       int_R_DATA_TEMPR69[1] ,int_R_DATA_TEMPR69[0] }), .DB_DETECT( int_DB_DETECT_NG[69] ), .SB_CORRECT(int_SB_CORRECT_NG[69] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[69] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[17] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[17] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_969 (.A(sel_R_DATA_TEMPR56[5] ), .B(sel_R_DATA_TEMPR57[5] ), .C(sel_R_DATA_TEMPR58[5] ), .D(sel_R_DATA_TEMPR59[5] ), .Y(OR4_969_Y));
    OR4 OR4_960 (.A(sel_R_DATA_TEMPR52[22] ), .B(sel_R_DATA_TEMPR53[22] ), 
        .C(sel_R_DATA_TEMPR54[22] ), .D(sel_R_DATA_TEMPR55[22] ), .Y(
        OR4_960_Y));
    OR4 OR4_197 (.A(sel_R_DATA_TEMPR4[3] ), .B(sel_R_DATA_TEMPR5[3] ), .C(sel_R_DATA_TEMPR6[3] ), .D(sel_R_DATA_TEMPR7[3] ), .Y(OR4_197_Y));
    OR4 OR4_1302 (.A(sel_R_DATA_TEMPR56[23] ), .B(sel_R_DATA_TEMPR57[23] ), 
        .C(sel_R_DATA_TEMPR58[23] ), .D(sel_R_DATA_TEMPR59[23] ), .Y(
        OR4_1302_Y));
    OR4 OR4_1149 (.A(sel_R_DATA_TEMPR44[26] ), .B(sel_R_DATA_TEMPR45[26] ), 
        .C(sel_R_DATA_TEMPR46[26] ), .D(sel_R_DATA_TEMPR47[26] ), .Y(
        OR4_1149_Y));
    OR4 OR4_1093 (.A(sel_R_DATA_TEMPR116[26] ), .B(sel_R_DATA_TEMPR117[26] ), 
        .C(sel_R_DATA_TEMPR118[26] ), .D(sel_R_DATA_TEMPR119[26] ), .Y(
        OR4_1093_Y));
    OR4 OR4_357 (.A(OR4_1347_Y), .B(OR4_815_Y), .C(OR4_1032_Y), .D(
        OR4_131_Y), .Y(OR4_357_Y));
    OR4 OR4_150 (.A(OR4_1369_Y), .B(OR4_1137_Y), .C(OR4_890_Y), .D(
        OR4_1109_Y), .Y(OR4_150_Y));
    OR4 OR4_434 (.A(sel_R_DATA_TEMPR104[3] ), .B(sel_R_DATA_TEMPR105[3] ), 
        .C(sel_R_DATA_TEMPR106[3] ), .D(sel_R_DATA_TEMPR107[3] ), .Y(
        OR4_434_Y));
    OR4 OR4_1202 (.A(\SB_CORRECT[36] ), .B(\SB_CORRECT[37] ), .C(
        \SB_CORRECT[38] ), .D(\SB_CORRECT[39] ), .Y(OR4_1202_Y));
    AND4 \AND4DB_DETECT[95]  (.A(sel_DB_DETECT_NG[95] ), .B(
        \BLKY2_pipe[23] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[95] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[26]  (.A(CFG3_14_Y), .B(
        CFG3_7_Y), .Y(\BLKX2[26] ));
    CFG3 #( .INIT(8'h20) )  CFG3_20 (.A(R_EN), .B(R_ADDR[15]), .C(
        R_ADDR[14]), .Y(CFG3_20_Y));
    OR4 OR4_163 (.A(OR4_406_Y), .B(OR4_885_Y), .C(OR4_175_Y), .D(
        OR4_395_Y), .Y(OR4_163_Y));
    OR4 OR4_1068 (.A(sel_R_DATA_TEMPR72[31] ), .B(sel_R_DATA_TEMPR73[31] ), 
        .C(sel_R_DATA_TEMPR74[31] ), .D(sel_R_DATA_TEMPR75[31] ), .Y(
        OR4_1068_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%38%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R38C0 (.A_DOUT({
        nc328, nc329, nc330, nc331, nc332,int_R_DATA_TEMPR38[31] , 
       int_R_DATA_TEMPR38[30] ,int_R_DATA_TEMPR38[29] , 
       int_R_DATA_TEMPR38[28] ,int_R_DATA_TEMPR38[27] , 
       int_R_DATA_TEMPR38[26] ,int_R_DATA_TEMPR38[25] , 
       int_R_DATA_TEMPR38[24] ,int_R_DATA_TEMPR38[23] , 
       int_R_DATA_TEMPR38[22] ,int_R_DATA_TEMPR38[21] , 
       int_R_DATA_TEMPR38[20] ,int_R_DATA_TEMPR38[19] , 
       int_R_DATA_TEMPR38[18] ,int_R_DATA_TEMPR38[17] }), .B_DOUT({nc333, 
        nc334, nc335,int_R_DATA_TEMPR38[16] ,int_R_DATA_TEMPR38[15] , 
       int_R_DATA_TEMPR38[14] ,int_R_DATA_TEMPR38[13] , 
       int_R_DATA_TEMPR38[12] ,int_R_DATA_TEMPR38[11] , 
       int_R_DATA_TEMPR38[10] ,int_R_DATA_TEMPR38[9] ,int_R_DATA_TEMPR38[8] , 
       int_R_DATA_TEMPR38[7] ,int_R_DATA_TEMPR38[6] ,int_R_DATA_TEMPR38[5] , 
       int_R_DATA_TEMPR38[4] ,int_R_DATA_TEMPR38[3] ,int_R_DATA_TEMPR38[2] , 
       int_R_DATA_TEMPR38[1] ,int_R_DATA_TEMPR38[0] }), .DB_DETECT( int_DB_DETECT_NG[38] ), .SB_CORRECT(int_SB_CORRECT_NG[38] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[38] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[9] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[9] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_758 (.A(OR4_1150_Y), .B(OR4_25_Y), .C(OR4_230_Y), .D(
        OR4_75_Y), .Y(OR4_758_Y));
    OR4 OR4_343 (.A(sel_R_DATA_TEMPR32[29] ), .B(sel_R_DATA_TEMPR33[29] ), 
        .C(sel_R_DATA_TEMPR34[29] ), .D(sel_R_DATA_TEMPR35[29] ), .Y(
        OR4_343_Y));
    OR4 OR4_740 (.A(sel_R_DATA_TEMPR124[3] ), .B(sel_R_DATA_TEMPR125[3] ), 
        .C(sel_R_DATA_TEMPR126[3] ), .D(sel_R_DATA_TEMPR127[3] ), .Y(
        OR4_740_Y));
    AND4 \AND4DB_DETECT[42]  (.A(sel_DB_DETECT_NG[42] ), .B(
        \BLKY2_pipe[10] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[42] ));
    DFN1E1 \DFN1E1BLKY2_pipe[15]  (.D(\BLKY2[15] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[15] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%35%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R35C0 (.A_DOUT({
        nc336, nc337, nc338, nc339, nc340,int_R_DATA_TEMPR35[31] , 
       int_R_DATA_TEMPR35[30] ,int_R_DATA_TEMPR35[29] , 
       int_R_DATA_TEMPR35[28] ,int_R_DATA_TEMPR35[27] , 
       int_R_DATA_TEMPR35[26] ,int_R_DATA_TEMPR35[25] , 
       int_R_DATA_TEMPR35[24] ,int_R_DATA_TEMPR35[23] , 
       int_R_DATA_TEMPR35[22] ,int_R_DATA_TEMPR35[21] , 
       int_R_DATA_TEMPR35[20] ,int_R_DATA_TEMPR35[19] , 
       int_R_DATA_TEMPR35[18] ,int_R_DATA_TEMPR35[17] }), .B_DOUT({nc341, 
        nc342, nc343,int_R_DATA_TEMPR35[16] ,int_R_DATA_TEMPR35[15] , 
       int_R_DATA_TEMPR35[14] ,int_R_DATA_TEMPR35[13] , 
       int_R_DATA_TEMPR35[12] ,int_R_DATA_TEMPR35[11] , 
       int_R_DATA_TEMPR35[10] ,int_R_DATA_TEMPR35[9] ,int_R_DATA_TEMPR35[8] , 
       int_R_DATA_TEMPR35[7] ,int_R_DATA_TEMPR35[6] ,int_R_DATA_TEMPR35[5] , 
       int_R_DATA_TEMPR35[4] ,int_R_DATA_TEMPR35[3] ,int_R_DATA_TEMPR35[2] , 
       int_R_DATA_TEMPR35[1] ,int_R_DATA_TEMPR35[0] }), .DB_DETECT( int_DB_DETECT_NG[35] ), .SB_CORRECT(int_SB_CORRECT_NG[35] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[35] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[8] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[8] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_336 (.A(sel_R_DATA_TEMPR112[5] ), .B(sel_R_DATA_TEMPR113[5] ), 
        .C(sel_R_DATA_TEMPR114[5] ), .D(sel_R_DATA_TEMPR115[5] ), .Y(
        OR4_336_Y));
    OR4 OR4_1280 (.A(sel_R_DATA_TEMPR4[19] ), .B(sel_R_DATA_TEMPR5[19] ), .C(sel_R_DATA_TEMPR6[19] ), .D(sel_R_DATA_TEMPR7[19] ), .Y(OR4_1280_Y));
    OR4 OR4_415 (.A(sel_R_DATA_TEMPR0[11] ), .B(sel_R_DATA_TEMPR1[11] ), .C(sel_R_DATA_TEMPR2[11] ), .D(sel_R_DATA_TEMPR3[11] ), .Y(OR4_415_Y));
    AND4 \AND4DB_DETECT[65]  (.A(sel_DB_DETECT_NG[65] ), .B(
        \BLKY2_pipe[16] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[65] ));
    OR4 OR4_793 (.A(\DB_DETECT[20] ), .B(\DB_DETECT[21] ), .C(
        \DB_DETECT[22] ), .D(\DB_DETECT[23] ), .Y(OR4_793_Y));
    OR4 OR4_442 (.A(sel_R_DATA_TEMPR112[17] ), .B(sel_R_DATA_TEMPR113[17] ), 
        .C(sel_R_DATA_TEMPR114[17] ), .D(sel_R_DATA_TEMPR115[17] ), .Y(
        OR4_442_Y));
    AND4 \AND4DB_DETECT[37]  (.A(sel_DB_DETECT_NG[37] ), .B(
        \BLKY2_pipe[9] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[37] ));
    OR4 OR4_1204 (.A(sel_R_DATA_TEMPR80[3] ), .B(sel_R_DATA_TEMPR81[3] ), .C(sel_R_DATA_TEMPR82[3] ), .D(sel_R_DATA_TEMPR83[3] ), .Y(OR4_1204_Y));
    OR4 OR4_294 (.A(OR4_1178_Y), .B(OR4_941_Y), .C(OR4_697_Y), .D(
        OR4_258_Y), .Y(OR4_294_Y));
    AND4 \AND4DB_DETECT[70]  (.A(sel_DB_DETECT_NG[70] ), .B(
        \BLKY2_pipe[17] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[70] ));
    OR4 OR4_449 (.A(OR4_714_Y), .B(OR4_218_Y), .C(OR4_662_Y), .D(
        OR4_1050_Y), .Y(OR4_449_Y));
    OR4 OR4_1174 (.A(sel_R_DATA_TEMPR32[27] ), .B(sel_R_DATA_TEMPR33[27] ), 
        .C(sel_R_DATA_TEMPR34[27] ), .D(sel_R_DATA_TEMPR35[27] ), .Y(
        OR4_1174_Y));
    OR4 OR4_505 (.A(sel_R_DATA_TEMPR0[23] ), .B(sel_R_DATA_TEMPR1[23] ), .C(sel_R_DATA_TEMPR2[23] ), .D(sel_R_DATA_TEMPR3[23] ), .Y(OR4_505_Y));
    OR4 OR4_1307 (.A(sel_R_DATA_TEMPR0[14] ), .B(sel_R_DATA_TEMPR1[14] ), .C(sel_R_DATA_TEMPR2[14] ), .D(sel_R_DATA_TEMPR3[14] ), .Y(OR4_1307_Y));
    OR4 \OR4_R_DATA[24]  (.A(OR4_1211_Y), .B(OR4_713_Y), .C(OR4_7_Y), 
        .D(OR4_602_Y), .Y(R_DATA[24]));
    OR4 OR4_85 (.A(sel_R_DATA_TEMPR24[11] ), .B(sel_R_DATA_TEMPR25[11] ), .C(sel_R_DATA_TEMPR26[11] ), .D(sel_R_DATA_TEMPR27[11] ), .Y(OR4_85_Y));
    OR4 OR4_1382 (.A(\DB_DETECT[36] ), .B(\DB_DETECT[37] ), .C(
        \DB_DETECT[38] ), .D(\DB_DETECT[39] ), .Y(OR4_1382_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[0]  (.D(\BLKY2[0] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[0] ));
    OR4 OR4_857 (.A(sel_R_DATA_TEMPR36[27] ), .B(sel_R_DATA_TEMPR37[27] ), 
        .C(sel_R_DATA_TEMPR38[27] ), .D(sel_R_DATA_TEMPR39[27] ), .Y(
        OR4_857_Y));
    AND4 \AND4DB_DETECT[83]  (.A(sel_DB_DETECT_NG[83] ), .B(
        \BLKY2_pipe[20] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[83] ));
    OR4 OR4_146 (.A(sel_R_DATA_TEMPR92[26] ), .B(sel_R_DATA_TEMPR93[26] ), 
        .C(sel_R_DATA_TEMPR94[26] ), .D(sel_R_DATA_TEMPR95[26] ), .Y(
        OR4_146_Y));
    OR4 OR4_158 (.A(sel_R_DATA_TEMPR12[18] ), .B(sel_R_DATA_TEMPR13[18] ), 
        .C(sel_R_DATA_TEMPR14[18] ), .D(sel_R_DATA_TEMPR15[18] ), .Y(
        OR4_158_Y));
    OR4 \OR4_R_DATA[12]  (.A(OR4_992_Y), .B(OR4_954_Y), .C(OR4_758_Y), 
        .D(OR4_140_Y), .Y(R_DATA[12]));
    OR4 OR4_954 (.A(OR4_372_Y), .B(OR4_108_Y), .C(OR4_97_Y), .D(
        OR4_751_Y), .Y(OR4_954_Y));
    OR4 OR4_1282 (.A(sel_R_DATA_TEMPR24[18] ), .B(sel_R_DATA_TEMPR25[18] ), 
        .C(sel_R_DATA_TEMPR26[18] ), .D(sel_R_DATA_TEMPR27[18] ), .Y(
        OR4_1282_Y));
    OR4 OR4_1146 (.A(OR4_336_Y), .B(OR4_554_Y), .C(OR4_709_Y), .D(
        OR4_1360_Y), .Y(OR4_1146_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_10 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_10_Y));
    OR4 OR4_581 (.A(sel_R_DATA_TEMPR32[15] ), .B(sel_R_DATA_TEMPR33[15] ), 
        .C(sel_R_DATA_TEMPR34[15] ), .D(sel_R_DATA_TEMPR35[15] ), .Y(
        OR4_581_Y));
    OR4 OR4_575 (.A(sel_R_DATA_TEMPR4[14] ), .B(sel_R_DATA_TEMPR5[14] ), .C(sel_R_DATA_TEMPR6[14] ), .D(sel_R_DATA_TEMPR7[14] ), .Y(OR4_575_Y));
    OR4 OR4_603 (.A(sel_R_DATA_TEMPR56[8] ), .B(sel_R_DATA_TEMPR57[8] ), .C(sel_R_DATA_TEMPR58[8] ), .D(sel_R_DATA_TEMPR59[8] ), .Y(OR4_603_Y));
    OR4 OR4_69 (.A(sel_R_DATA_TEMPR116[22] ), .B(sel_R_DATA_TEMPR117[22] ), 
        .C(sel_R_DATA_TEMPR118[22] ), .D(sel_R_DATA_TEMPR119[22] ), .Y(
        OR4_69_Y));
    OR4 OR4_1241 (.A(OR4_581_Y), .B(OR4_124_Y), .C(OR4_104_Y), .D(
        OR4_764_Y), .Y(OR4_1241_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%16%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R16C0 (.A_DOUT({
        nc344, nc345, nc346, nc347, nc348,int_R_DATA_TEMPR16[31] , 
       int_R_DATA_TEMPR16[30] ,int_R_DATA_TEMPR16[29] , 
       int_R_DATA_TEMPR16[28] ,int_R_DATA_TEMPR16[27] , 
       int_R_DATA_TEMPR16[26] ,int_R_DATA_TEMPR16[25] , 
       int_R_DATA_TEMPR16[24] ,int_R_DATA_TEMPR16[23] , 
       int_R_DATA_TEMPR16[22] ,int_R_DATA_TEMPR16[21] , 
       int_R_DATA_TEMPR16[20] ,int_R_DATA_TEMPR16[19] , 
       int_R_DATA_TEMPR16[18] ,int_R_DATA_TEMPR16[17] }), .B_DOUT({nc349, 
        nc350, nc351,int_R_DATA_TEMPR16[16] ,int_R_DATA_TEMPR16[15] , 
       int_R_DATA_TEMPR16[14] ,int_R_DATA_TEMPR16[13] , 
       int_R_DATA_TEMPR16[12] ,int_R_DATA_TEMPR16[11] , 
       int_R_DATA_TEMPR16[10] ,int_R_DATA_TEMPR16[9] ,int_R_DATA_TEMPR16[8] , 
       int_R_DATA_TEMPR16[7] ,int_R_DATA_TEMPR16[6] ,int_R_DATA_TEMPR16[5] , 
       int_R_DATA_TEMPR16[4] ,int_R_DATA_TEMPR16[3] ,int_R_DATA_TEMPR16[2] , 
       int_R_DATA_TEMPR16[1] ,int_R_DATA_TEMPR16[0] }), .DB_DETECT( int_DB_DETECT_NG[16] ), .SB_CORRECT(int_SB_CORRECT_NG[16] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[16] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[4] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1148 (.A(OR4_792_Y), .B(OR2_0_Y), .C(sel_R_DATA_TEMPR86[16] ), 
        .D(sel_R_DATA_TEMPR87[16] ), .Y(OR4_1148_Y));
    OR4 OR4_1157 (.A(sel_R_DATA_TEMPR24[25] ), .B(sel_R_DATA_TEMPR25[25] ), 
        .C(sel_R_DATA_TEMPR26[25] ), .D(sel_R_DATA_TEMPR27[25] ), .Y(
        OR4_1157_Y));
    OR4 OR4_227 (.A(sel_R_DATA_TEMPR120[1] ), .B(sel_R_DATA_TEMPR121[1] ), 
        .C(sel_R_DATA_TEMPR122[1] ), .D(sel_R_DATA_TEMPR123[1] ), .Y(
        OR4_227_Y));
    OR4 OR4_1278 (.A(sel_R_DATA_TEMPR76[26] ), .B(sel_R_DATA_TEMPR77[26] ), 
        .C(sel_R_DATA_TEMPR78[26] ), .D(sel_R_DATA_TEMPR79[26] ), .Y(
        OR4_1278_Y));
    OR4 OR4_673 (.A(sel_R_DATA_TEMPR24[26] ), .B(sel_R_DATA_TEMPR25[26] ), 
        .C(sel_R_DATA_TEMPR26[26] ), .D(sel_R_DATA_TEMPR27[26] ), .Y(
        OR4_673_Y));
    OR4 OR4_1217 (.A(OR4_228_Y), .B(OR4_942_Y), .C(OR4_21_Y), .D(
        OR4_887_Y), .Y(OR4_1217_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[21]  (.A(CFG3_11_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[21] ));
    OR4 OR4_395 (.A(sel_R_DATA_TEMPR60[20] ), .B(sel_R_DATA_TEMPR61[20] ), 
        .C(sel_R_DATA_TEMPR62[20] ), .D(sel_R_DATA_TEMPR63[20] ), .Y(
        OR4_395_Y));
    OR4 OR4_414 (.A(sel_R_DATA_TEMPR60[11] ), .B(sel_R_DATA_TEMPR61[11] ), 
        .C(sel_R_DATA_TEMPR62[11] ), .D(sel_R_DATA_TEMPR63[11] ), .Y(
        OR4_414_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[19]  (.D(\BLKY2[19] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[19] ));
    OR4 OR4_127 (.A(sel_R_DATA_TEMPR60[23] ), .B(sel_R_DATA_TEMPR61[23] ), 
        .C(sel_R_DATA_TEMPR62[23] ), .D(sel_R_DATA_TEMPR63[23] ), .Y(
        OR4_127_Y));
    OR4 OR4_1284 (.A(sel_R_DATA_TEMPR96[10] ), .B(sel_R_DATA_TEMPR97[10] ), 
        .C(sel_R_DATA_TEMPR98[10] ), .D(sel_R_DATA_TEMPR99[10] ), .Y(
        OR4_1284_Y));
    OR4 OR4_860 (.A(sel_R_DATA_TEMPR104[21] ), .B(sel_R_DATA_TEMPR105[21] ), 
        .C(sel_R_DATA_TEMPR106[21] ), .D(sel_R_DATA_TEMPR107[21] ), .Y(
        OR4_860_Y));
    OR4 OR4_348 (.A(sel_R_DATA_TEMPR80[26] ), .B(sel_R_DATA_TEMPR81[26] ), 
        .C(sel_R_DATA_TEMPR82[26] ), .D(sel_R_DATA_TEMPR83[26] ), .Y(
        OR4_348_Y));
    OR4 OR4_1098 (.A(sel_R_DATA_TEMPR108[16] ), .B(sel_R_DATA_TEMPR109[16] ), 
        .C(sel_R_DATA_TEMPR110[16] ), .D(sel_R_DATA_TEMPR111[16] ), .Y(
        OR4_1098_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%82%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R82C0 (.A_DOUT({
        nc352, nc353, nc354, nc355, nc356,int_R_DATA_TEMPR82[31] , 
       int_R_DATA_TEMPR82[30] ,int_R_DATA_TEMPR82[29] , 
       int_R_DATA_TEMPR82[28] ,int_R_DATA_TEMPR82[27] , 
       int_R_DATA_TEMPR82[26] ,int_R_DATA_TEMPR82[25] , 
       int_R_DATA_TEMPR82[24] ,int_R_DATA_TEMPR82[23] , 
       int_R_DATA_TEMPR82[22] ,int_R_DATA_TEMPR82[21] , 
       int_R_DATA_TEMPR82[20] ,int_R_DATA_TEMPR82[19] , 
       int_R_DATA_TEMPR82[18] ,int_R_DATA_TEMPR82[17] }), .B_DOUT({nc357, 
        nc358, nc359,int_R_DATA_TEMPR82[16] ,int_R_DATA_TEMPR82[15] , 
       int_R_DATA_TEMPR82[14] ,int_R_DATA_TEMPR82[13] , 
       int_R_DATA_TEMPR82[12] ,int_R_DATA_TEMPR82[11] , 
       int_R_DATA_TEMPR82[10] ,int_R_DATA_TEMPR82[9] ,int_R_DATA_TEMPR82[8] , 
       int_R_DATA_TEMPR82[7] ,int_R_DATA_TEMPR82[6] ,int_R_DATA_TEMPR82[5] , 
       int_R_DATA_TEMPR82[4] ,int_R_DATA_TEMPR82[3] ,int_R_DATA_TEMPR82[2] , 
       int_R_DATA_TEMPR82[1] ,int_R_DATA_TEMPR82[0] }), .DB_DETECT( int_DB_DETECT_NG[82] ), .SB_CORRECT(int_SB_CORRECT_NG[82] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[82] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[20] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[20] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_162 (.A(OR4_483_Y), .B(OR4_960_Y), .C(OR4_259_Y), .D(
        OR4_476_Y), .Y(OR4_162_Y));
    OR4 OR4_1387 (.A(sel_R_DATA_TEMPR36[23] ), .B(sel_R_DATA_TEMPR37[23] ), 
        .C(sel_R_DATA_TEMPR38[23] ), .D(sel_R_DATA_TEMPR39[23] ), .Y(
        OR4_1387_Y));
    OR4 OR4_282 (.A(sel_R_DATA_TEMPR40[26] ), .B(sel_R_DATA_TEMPR41[26] ), 
        .C(sel_R_DATA_TEMPR42[26] ), .D(sel_R_DATA_TEMPR43[26] ), .Y(
        OR4_282_Y));
    OR4 OR4_965 (.A(sel_R_DATA_TEMPR40[18] ), .B(sel_R_DATA_TEMPR41[18] ), 
        .C(sel_R_DATA_TEMPR42[18] ), .D(sel_R_DATA_TEMPR43[18] ), .Y(
        OR4_965_Y));
    OR4 OR4_316 (.A(sel_R_DATA_TEMPR60[5] ), .B(sel_R_DATA_TEMPR61[5] ), .C(sel_R_DATA_TEMPR62[5] ), .D(sel_R_DATA_TEMPR63[5] ), .Y(OR4_316_Y));
    OR4 OR4_1314 (.A(sel_R_DATA_TEMPR120[15] ), .B(sel_R_DATA_TEMPR121[15] ), 
        .C(sel_R_DATA_TEMPR122[15] ), .D(sel_R_DATA_TEMPR123[15] ), .Y(
        OR4_1314_Y));
    OR4 OR4_909 (.A(sel_R_DATA_TEMPR64[9] ), .B(sel_R_DATA_TEMPR65[9] ), .C(sel_R_DATA_TEMPR66[9] ), .D(sel_R_DATA_TEMPR67[9] ), .Y(OR4_909_Y));
    OR4 OR4_900 (.A(sel_R_DATA_TEMPR104[17] ), .B(sel_R_DATA_TEMPR105[17] ), 
        .C(sel_R_DATA_TEMPR106[17] ), .D(sel_R_DATA_TEMPR107[17] ), .Y(
        OR4_900_Y));
    OR4 OR4_134 (.A(OR4_358_Y), .B(OR4_839_Y), .C(OR4_120_Y), .D(
        OR4_349_Y), .Y(OR4_134_Y));
    OR4 OR4_723 (.A(OR4_1198_Y), .B(OR4_904_Y), .C(OR4_881_Y), .D(
        OR4_356_Y), .Y(OR4_723_Y));
    OR4 OR4_979 (.A(sel_R_DATA_TEMPR36[29] ), .B(sel_R_DATA_TEMPR37[29] ), 
        .C(sel_R_DATA_TEMPR38[29] ), .D(sel_R_DATA_TEMPR39[29] ), .Y(
        OR4_979_Y));
    OR4 OR4_970 (.A(sel_R_DATA_TEMPR56[7] ), .B(sel_R_DATA_TEMPR57[7] ), .C(sel_R_DATA_TEMPR58[7] ), .D(sel_R_DATA_TEMPR59[7] ), .Y(OR4_970_Y));
    OR4 OR4_1067 (.A(OR4_1114_Y), .B(OR4_877_Y), .C(OR4_640_Y), .D(
        OR4_1076_Y), .Y(OR4_1067_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%109%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R109C0 (.A_DOUT({
        nc360, nc361, nc362, nc363, nc364,int_R_DATA_TEMPR109[31] , 
       int_R_DATA_TEMPR109[30] ,int_R_DATA_TEMPR109[29] , 
       int_R_DATA_TEMPR109[28] ,int_R_DATA_TEMPR109[27] , 
       int_R_DATA_TEMPR109[26] ,int_R_DATA_TEMPR109[25] , 
       int_R_DATA_TEMPR109[24] ,int_R_DATA_TEMPR109[23] , 
       int_R_DATA_TEMPR109[22] ,int_R_DATA_TEMPR109[21] , 
       int_R_DATA_TEMPR109[20] ,int_R_DATA_TEMPR109[19] , 
       int_R_DATA_TEMPR109[18] ,int_R_DATA_TEMPR109[17] }), .B_DOUT({nc365, 
        nc366, nc367,int_R_DATA_TEMPR109[16] ,int_R_DATA_TEMPR109[15] , 
       int_R_DATA_TEMPR109[14] ,int_R_DATA_TEMPR109[13] , 
       int_R_DATA_TEMPR109[12] ,int_R_DATA_TEMPR109[11] , 
       int_R_DATA_TEMPR109[10] ,int_R_DATA_TEMPR109[9] , 
       int_R_DATA_TEMPR109[8] ,int_R_DATA_TEMPR109[7] , 
       int_R_DATA_TEMPR109[6] ,int_R_DATA_TEMPR109[5] , 
       int_R_DATA_TEMPR109[4] ,int_R_DATA_TEMPR109[3] , 
       int_R_DATA_TEMPR109[2] ,int_R_DATA_TEMPR109[1] , 
       int_R_DATA_TEMPR109[0] }), .DB_DETECT(int_DB_DETECT_NG[109] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[109] ), .ACCESS_BUSY(
        ACCESS_BUSY[109] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[27] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[27] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_103 (.A(sel_R_DATA_TEMPR48[11] ), .B(sel_R_DATA_TEMPR49[11] ), 
        .C(sel_R_DATA_TEMPR50[11] ), .D(sel_R_DATA_TEMPR51[11] ), .Y(
        OR4_103_Y));
    AND4 \AND4SB_CORRECT[25]  (.A(sel_SB_CORRECT_NG[25] ), .B(
        \BLKY2_pipe[6] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[25] ));
    AND4 \AND4SB_CORRECT[26]  (.A(sel_SB_CORRECT_NG[26] ), .B(
        \BLKY2_pipe[6] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[26] ));
    OR4 OR4_224 (.A(sel_R_DATA_TEMPR88[10] ), .B(sel_R_DATA_TEMPR89[10] ), 
        .C(sel_R_DATA_TEMPR90[10] ), .D(sel_R_DATA_TEMPR91[10] ), .Y(
        OR4_224_Y));
    DFN1E1 \DFN1E1BLKY1_pipe[1]  (.D(R_ADDR[10]), .CLK(CLK), .E(VCC), 
        .Q(\BLKY1_pipe[1] ));
    OR4 OR4_149 (.A(sel_R_DATA_TEMPR96[29] ), .B(sel_R_DATA_TEMPR97[29] ), 
        .C(sel_R_DATA_TEMPR98[29] ), .D(sel_R_DATA_TEMPR99[29] ), .Y(
        OR4_149_Y));
    OR4 OR4_792 (.A(sel_R_DATA_TEMPR80[16] ), .B(sel_R_DATA_TEMPR81[16] ), 
        .C(sel_R_DATA_TEMPR82[16] ), .D(sel_R_DATA_TEMPR83[16] ), .Y(
        OR4_792_Y));
    AND4 \AND4DB_DETECT[3]  (.A(sel_DB_DETECT_NG[3] ), .B(
        \BLKY2_pipe[0] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[3] ));
    OR4 OR4_380 (.A(sel_R_DATA_TEMPR68[6] ), .B(sel_R_DATA_TEMPR69[6] ), .C(sel_R_DATA_TEMPR70[6] ), .D(sel_R_DATA_TEMPR71[6] ), .Y(OR4_380_Y));
    OR4 OR4_933 (.A(sel_R_DATA_TEMPR20[15] ), .B(sel_R_DATA_TEMPR21[15] ), 
        .C(sel_R_DATA_TEMPR22[15] ), .D(sel_R_DATA_TEMPR23[15] ), .Y(
        OR4_933_Y));
    OR4 \OR4_R_DATA[13]  (.A(OR4_832_Y), .B(OR4_486_Y), .C(OR4_435_Y), 
        .D(OR4_388_Y), .Y(R_DATA[13]));
    OR4 OR4_173 (.A(sel_R_DATA_TEMPR92[8] ), .B(sel_R_DATA_TEMPR93[8] ), .C(sel_R_DATA_TEMPR94[8] ), .D(sel_R_DATA_TEMPR95[8] ), .Y(OR4_173_Y));
    OR4 OR4_269 (.A(sel_R_DATA_TEMPR28[5] ), .B(sel_R_DATA_TEMPR29[5] ), .C(sel_R_DATA_TEMPR30[5] ), .D(sel_R_DATA_TEMPR31[5] ), .Y(OR4_269_Y));
    OR4 OR4_996 (.A(sel_R_DATA_TEMPR72[8] ), .B(sel_R_DATA_TEMPR73[8] ), .C(sel_R_DATA_TEMPR74[8] ), .D(sel_R_DATA_TEMPR75[8] ), .Y(OR4_996_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[31]  (.A(CFG3_23_Y), .B(
        CFG3_7_Y), .Y(\BLKX2[31] ));
    OR4 OR4_836 (.A(sel_R_DATA_TEMPR96[20] ), .B(sel_R_DATA_TEMPR97[20] ), 
        .C(sel_R_DATA_TEMPR98[20] ), .D(sel_R_DATA_TEMPR99[20] ), .Y(
        OR4_836_Y));
    AND4 \AND4SB_CORRECT[79]  (.A(sel_SB_CORRECT_NG[79] ), .B(
        \BLKY2_pipe[19] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[79] ));
    OR4 OR4_731 (.A(OR4_179_Y), .B(OR4_41_Y), .C(OR4_144_Y), .D(
        OR4_309_Y), .Y(OR4_731_Y));
    OR4 OR4_695 (.A(sel_R_DATA_TEMPR48[31] ), .B(sel_R_DATA_TEMPR49[31] ), 
        .C(sel_R_DATA_TEMPR50[31] ), .D(sel_R_DATA_TEMPR51[31] ), .Y(
        OR4_695_Y));
    OR4 OR4_62 (.A(sel_R_DATA_TEMPR36[28] ), .B(sel_R_DATA_TEMPR37[28] ), .C(sel_R_DATA_TEMPR38[28] ), .D(sel_R_DATA_TEMPR39[28] ), .Y(OR4_62_Y));
    OR4 OR4_883 (.A(sel_R_DATA_TEMPR12[15] ), .B(sel_R_DATA_TEMPR13[15] ), 
        .C(sel_R_DATA_TEMPR14[15] ), .D(sel_R_DATA_TEMPR15[15] ), .Y(
        OR4_883_Y));
    AND4 \AND4DB_DETECT[104]  (.A(sel_DB_DETECT_NG[104] ), .B(
        \BLKY2_pipe[26] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[104] ));
    OR4 OR4_1175 (.A(sel_R_DATA_TEMPR80[18] ), .B(sel_R_DATA_TEMPR81[18] ), 
        .C(sel_R_DATA_TEMPR82[18] ), .D(sel_R_DATA_TEMPR83[18] ), .Y(
        OR4_1175_Y));
    OR4 OR4_941 (.A(sel_R_DATA_TEMPR68[28] ), .B(sel_R_DATA_TEMPR69[28] ), 
        .C(sel_R_DATA_TEMPR70[28] ), .D(sel_R_DATA_TEMPR71[28] ), .Y(
        OR4_941_Y));
    OR4 OR4_1319 (.A(OR4_221_Y), .B(OR4_263_Y), .C(OR4_700_Y), .D(
        OR4_1087_Y), .Y(OR4_1319_Y));
    OR4 OR4_38 (.A(sel_R_DATA_TEMPR120[14] ), .B(sel_R_DATA_TEMPR121[14] ), 
        .C(sel_R_DATA_TEMPR122[14] ), .D(sel_R_DATA_TEMPR123[14] ), .Y(
        OR4_38_Y));
    OR4 OR4_1250 (.A(OR4_76_Y), .B(OR2_23_Y), .C(sel_R_DATA_TEMPR86[27] ), 
        .D(sel_R_DATA_TEMPR87[27] ), .Y(OR4_1250_Y));
    OR4 OR4_1071 (.A(sel_R_DATA_TEMPR116[31] ), .B(sel_R_DATA_TEMPR117[31] ), 
        .C(sel_R_DATA_TEMPR118[31] ), .D(sel_R_DATA_TEMPR119[31] ), .Y(
        OR4_1071_Y));
    OR4 OR4_1010 (.A(OR4_899_Y), .B(OR4_606_Y), .C(OR4_919_Y), .D(
        OR4_163_Y), .Y(OR4_1010_Y));
    AND4 \AND4SB_CORRECT[82]  (.A(sel_SB_CORRECT_NG[82] ), .B(
        \BLKY2_pipe[20] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[82] ));
    OR4 OR4_325 (.A(OR4_867_Y), .B(OR4_1351_Y), .C(OR4_552_Y), .D(
        OR4_1120_Y), .Y(OR4_325_Y));
    DFN1E1 \DFN1E1BLKY0_pipe[0]  (.D(\BLKY0[0] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY0_pipe[0] ));
    OR4 OR4_1306 (.A(\DB_DETECT[68] ), .B(\DB_DETECT[69] ), .C(
        \DB_DETECT[70] ), .D(\DB_DETECT[71] ), .Y(OR4_1306_Y));
    OR4 OR4_536 (.A(sel_R_DATA_TEMPR56[4] ), .B(sel_R_DATA_TEMPR57[4] ), .C(sel_R_DATA_TEMPR58[4] ), .D(sel_R_DATA_TEMPR59[4] ), .Y(OR4_536_Y));
    OR4 OR4_869 (.A(OR4_1118_Y), .B(OR4_1383_Y), .C(OR4_896_Y), .D(
        OR4_248_Y), .Y(OR4_869_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%126%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R126C0 (.A_DOUT({
        nc368, nc369, nc370, nc371, nc372,int_R_DATA_TEMPR126[31] , 
       int_R_DATA_TEMPR126[30] ,int_R_DATA_TEMPR126[29] , 
       int_R_DATA_TEMPR126[28] ,int_R_DATA_TEMPR126[27] , 
       int_R_DATA_TEMPR126[26] ,int_R_DATA_TEMPR126[25] , 
       int_R_DATA_TEMPR126[24] ,int_R_DATA_TEMPR126[23] , 
       int_R_DATA_TEMPR126[22] ,int_R_DATA_TEMPR126[21] , 
       int_R_DATA_TEMPR126[20] ,int_R_DATA_TEMPR126[19] , 
       int_R_DATA_TEMPR126[18] ,int_R_DATA_TEMPR126[17] }), .B_DOUT({nc373, 
        nc374, nc375,int_R_DATA_TEMPR126[16] ,int_R_DATA_TEMPR126[15] , 
       int_R_DATA_TEMPR126[14] ,int_R_DATA_TEMPR126[13] , 
       int_R_DATA_TEMPR126[12] ,int_R_DATA_TEMPR126[11] , 
       int_R_DATA_TEMPR126[10] ,int_R_DATA_TEMPR126[9] , 
       int_R_DATA_TEMPR126[8] ,int_R_DATA_TEMPR126[7] , 
       int_R_DATA_TEMPR126[6] ,int_R_DATA_TEMPR126[5] , 
       int_R_DATA_TEMPR126[4] ,int_R_DATA_TEMPR126[3] , 
       int_R_DATA_TEMPR126[2] ,int_R_DATA_TEMPR126[1] , 
       int_R_DATA_TEMPR126[0] }), .DB_DETECT(int_DB_DETECT_NG[126] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[126] ), .ACCESS_BUSY(
        ACCESS_BUSY[126] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[31] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[31] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1352 (.A(sel_R_DATA_TEMPR32[28] ), .B(sel_R_DATA_TEMPR33[28] ), 
        .C(sel_R_DATA_TEMPR34[28] ), .D(sel_R_DATA_TEMPR35[28] ), .Y(
        OR4_1352_Y));
    AND4 \AND4SB_CORRECT[65]  (.A(sel_SB_CORRECT_NG[65] ), .B(
        \BLKY2_pipe[16] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[65] ));
    AND4 \AND4SB_CORRECT[66]  (.A(sel_SB_CORRECT_NG[66] ), .B(
        \BLKY2_pipe[16] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[66] ));
    OR4 OR4_114 (.A(sel_R_DATA_TEMPR20[2] ), .B(sel_R_DATA_TEMPR21[2] ), .C(sel_R_DATA_TEMPR22[2] ), .D(sel_R_DATA_TEMPR23[2] ), .Y(OR4_114_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[28]  (.D(\BLKY2[28] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[28] ));
    OR4 OR4_155 (.A(\SB_CORRECT[12] ), .B(\SB_CORRECT[13] ), .C(
        \SB_CORRECT[14] ), .D(\SB_CORRECT[15] ), .Y(OR4_155_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[6]  (.A(CFG3_10_Y), .B(
        CFG3_12_Y), .Y(\BLKX2[6] ));
    OR4 OR4_1252 (.A(sel_R_DATA_TEMPR88[2] ), .B(sel_R_DATA_TEMPR89[2] ), .C(sel_R_DATA_TEMPR90[2] ), .D(sel_R_DATA_TEMPR91[2] ), .Y(OR4_1252_Y));
    OR4 OR4_800 (.A(OR4_1332_Y), .B(OR4_202_Y), .C(OR4_1008_Y), .D(
        OR4_846_Y), .Y(OR4_800_Y));
    AND4 \AND4DB_DETECT[114]  (.A(sel_DB_DETECT_NG[114] ), .B(
        \BLKY2_pipe[28] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[114] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%78%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R78C0 (.A_DOUT({
        nc376, nc377, nc378, nc379, nc380,int_R_DATA_TEMPR78[31] , 
       int_R_DATA_TEMPR78[30] ,int_R_DATA_TEMPR78[29] , 
       int_R_DATA_TEMPR78[28] ,int_R_DATA_TEMPR78[27] , 
       int_R_DATA_TEMPR78[26] ,int_R_DATA_TEMPR78[25] , 
       int_R_DATA_TEMPR78[24] ,int_R_DATA_TEMPR78[23] , 
       int_R_DATA_TEMPR78[22] ,int_R_DATA_TEMPR78[21] , 
       int_R_DATA_TEMPR78[20] ,int_R_DATA_TEMPR78[19] , 
       int_R_DATA_TEMPR78[18] ,int_R_DATA_TEMPR78[17] }), .B_DOUT({nc381, 
        nc382, nc383,int_R_DATA_TEMPR78[16] ,int_R_DATA_TEMPR78[15] , 
       int_R_DATA_TEMPR78[14] ,int_R_DATA_TEMPR78[13] , 
       int_R_DATA_TEMPR78[12] ,int_R_DATA_TEMPR78[11] , 
       int_R_DATA_TEMPR78[10] ,int_R_DATA_TEMPR78[9] ,int_R_DATA_TEMPR78[8] , 
       int_R_DATA_TEMPR78[7] ,int_R_DATA_TEMPR78[6] ,int_R_DATA_TEMPR78[5] , 
       int_R_DATA_TEMPR78[4] ,int_R_DATA_TEMPR78[3] ,int_R_DATA_TEMPR78[2] , 
       int_R_DATA_TEMPR78[1] ,int_R_DATA_TEMPR78[0] }), .DB_DETECT( int_DB_DETECT_NG[78] ), .SB_CORRECT(int_SB_CORRECT_NG[78] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[78] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[19] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[19] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1097 (.A(sel_R_DATA_TEMPR44[11] ), .B(sel_R_DATA_TEMPR45[11] ), 
        .C(sel_R_DATA_TEMPR46[11] ), .D(sel_R_DATA_TEMPR47[11] ), .Y(
        OR4_1097_Y));
    OR4 OR4_1073 (.A(sel_R_DATA_TEMPR52[8] ), .B(sel_R_DATA_TEMPR53[8] ), .C(sel_R_DATA_TEMPR54[8] ), .D(sel_R_DATA_TEMPR55[8] ), .Y(OR4_1073_Y));
    AND4 \AND4SB_CORRECT[33]  (.A(sel_SB_CORRECT_NG[33] ), .B(
        \BLKY2_pipe[8] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[33] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[14]  (.A(CFG3_10_Y), .B(
        CFG3_4_Y), .Y(\BLKX2[14] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%59%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R59C0 (.A_DOUT({
        nc384, nc385, nc386, nc387, nc388,int_R_DATA_TEMPR59[31] , 
       int_R_DATA_TEMPR59[30] ,int_R_DATA_TEMPR59[29] , 
       int_R_DATA_TEMPR59[28] ,int_R_DATA_TEMPR59[27] , 
       int_R_DATA_TEMPR59[26] ,int_R_DATA_TEMPR59[25] , 
       int_R_DATA_TEMPR59[24] ,int_R_DATA_TEMPR59[23] , 
       int_R_DATA_TEMPR59[22] ,int_R_DATA_TEMPR59[21] , 
       int_R_DATA_TEMPR59[20] ,int_R_DATA_TEMPR59[19] , 
       int_R_DATA_TEMPR59[18] ,int_R_DATA_TEMPR59[17] }), .B_DOUT({nc389, 
        nc390, nc391,int_R_DATA_TEMPR59[16] ,int_R_DATA_TEMPR59[15] , 
       int_R_DATA_TEMPR59[14] ,int_R_DATA_TEMPR59[13] , 
       int_R_DATA_TEMPR59[12] ,int_R_DATA_TEMPR59[11] , 
       int_R_DATA_TEMPR59[10] ,int_R_DATA_TEMPR59[9] ,int_R_DATA_TEMPR59[8] , 
       int_R_DATA_TEMPR59[7] ,int_R_DATA_TEMPR59[6] ,int_R_DATA_TEMPR59[5] , 
       int_R_DATA_TEMPR59[4] ,int_R_DATA_TEMPR59[3] ,int_R_DATA_TEMPR59[2] , 
       int_R_DATA_TEMPR59[1] ,int_R_DATA_TEMPR59[0] }), .DB_DETECT( int_DB_DETECT_NG[59] ), .SB_CORRECT(int_SB_CORRECT_NG[59] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[59] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[14] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[14] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%75%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R75C0 (.A_DOUT({
        nc392, nc393, nc394, nc395, nc396,int_R_DATA_TEMPR75[31] , 
       int_R_DATA_TEMPR75[30] ,int_R_DATA_TEMPR75[29] , 
       int_R_DATA_TEMPR75[28] ,int_R_DATA_TEMPR75[27] , 
       int_R_DATA_TEMPR75[26] ,int_R_DATA_TEMPR75[25] , 
       int_R_DATA_TEMPR75[24] ,int_R_DATA_TEMPR75[23] , 
       int_R_DATA_TEMPR75[22] ,int_R_DATA_TEMPR75[21] , 
       int_R_DATA_TEMPR75[20] ,int_R_DATA_TEMPR75[19] , 
       int_R_DATA_TEMPR75[18] ,int_R_DATA_TEMPR75[17] }), .B_DOUT({nc397, 
        nc398, nc399,int_R_DATA_TEMPR75[16] ,int_R_DATA_TEMPR75[15] , 
       int_R_DATA_TEMPR75[14] ,int_R_DATA_TEMPR75[13] , 
       int_R_DATA_TEMPR75[12] ,int_R_DATA_TEMPR75[11] , 
       int_R_DATA_TEMPR75[10] ,int_R_DATA_TEMPR75[9] ,int_R_DATA_TEMPR75[8] , 
       int_R_DATA_TEMPR75[7] ,int_R_DATA_TEMPR75[6] ,int_R_DATA_TEMPR75[5] , 
       int_R_DATA_TEMPR75[4] ,int_R_DATA_TEMPR75[3] ,int_R_DATA_TEMPR75[2] , 
       int_R_DATA_TEMPR75[1] ,int_R_DATA_TEMPR75[0] }), .DB_DETECT( int_DB_DETECT_NG[75] ), .SB_CORRECT(int_SB_CORRECT_NG[75] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[75] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[18] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[18] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_457 (.A(sel_R_DATA_TEMPR4[30] ), .B(sel_R_DATA_TEMPR5[30] ), .C(sel_R_DATA_TEMPR6[30] ), .D(sel_R_DATA_TEMPR7[30] ), .Y(OR4_457_Y));
    OR4 OR4_102 (.A(\SB_CORRECT[8] ), .B(\SB_CORRECT[9] ), .C(
        \SB_CORRECT[10] ), .D(\SB_CORRECT[11] ), .Y(OR4_102_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[25]  (.A(CFG3_15_Y), .B(
        CFG3_3_Y), .Y(\BLKY2[25] ));
    OR4 OR4_905 (.A(sel_R_DATA_TEMPR48[3] ), .B(sel_R_DATA_TEMPR49[3] ), .C(sel_R_DATA_TEMPR50[3] ), .D(sel_R_DATA_TEMPR51[3] ), .Y(OR4_905_Y));
    OR4 OR4_870 (.A(sel_R_DATA_TEMPR60[13] ), .B(sel_R_DATA_TEMPR61[13] ), 
        .C(sel_R_DATA_TEMPR62[13] ), .D(sel_R_DATA_TEMPR63[13] ), .Y(
        OR4_870_Y));
    AND4 \AND4DB_DETECT[125]  (.A(sel_DB_DETECT_NG[125] ), .B(
        \BLKY2_pipe[31] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[125] ));
    INV \INVBLKY0[0]  (.A(R_ADDR[9]), .Y(\BLKY0[0] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%67%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R67C0 (.A_DOUT({
        nc400, nc401, nc402, nc403, nc404,int_R_DATA_TEMPR67[31] , 
       int_R_DATA_TEMPR67[30] ,int_R_DATA_TEMPR67[29] , 
       int_R_DATA_TEMPR67[28] ,int_R_DATA_TEMPR67[27] , 
       int_R_DATA_TEMPR67[26] ,int_R_DATA_TEMPR67[25] , 
       int_R_DATA_TEMPR67[24] ,int_R_DATA_TEMPR67[23] , 
       int_R_DATA_TEMPR67[22] ,int_R_DATA_TEMPR67[21] , 
       int_R_DATA_TEMPR67[20] ,int_R_DATA_TEMPR67[19] , 
       int_R_DATA_TEMPR67[18] ,int_R_DATA_TEMPR67[17] }), .B_DOUT({nc405, 
        nc406, nc407,int_R_DATA_TEMPR67[16] ,int_R_DATA_TEMPR67[15] , 
       int_R_DATA_TEMPR67[14] ,int_R_DATA_TEMPR67[13] , 
       int_R_DATA_TEMPR67[12] ,int_R_DATA_TEMPR67[11] , 
       int_R_DATA_TEMPR67[10] ,int_R_DATA_TEMPR67[9] ,int_R_DATA_TEMPR67[8] , 
       int_R_DATA_TEMPR67[7] ,int_R_DATA_TEMPR67[6] ,int_R_DATA_TEMPR67[5] , 
       int_R_DATA_TEMPR67[4] ,int_R_DATA_TEMPR67[3] ,int_R_DATA_TEMPR67[2] , 
       int_R_DATA_TEMPR67[1] ,int_R_DATA_TEMPR67[0] }), .DB_DETECT( int_DB_DETECT_NG[67] ), .SB_CORRECT(int_SB_CORRECT_NG[67] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[67] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[16] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[16] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_913 (.A(OR4_141_Y), .B(OR4_6_Y), .C(OR4_107_Y), .D(
        OR4_445_Y), .Y(OR4_913_Y));
    OR4 OR4_690 (.A(sel_R_DATA_TEMPR52[28] ), .B(sel_R_DATA_TEMPR53[28] ), 
        .C(sel_R_DATA_TEMPR54[28] ), .D(sel_R_DATA_TEMPR55[28] ), .Y(
        OR4_690_Y));
    OR4 OR4_1133 (.A(sel_R_DATA_TEMPR116[10] ), .B(sel_R_DATA_TEMPR117[10] ), 
        .C(sel_R_DATA_TEMPR118[10] ), .D(sel_R_DATA_TEMPR119[10] ), .Y(
        OR4_1133_Y));
    OR4 OR4_722 (.A(OR4_669_Y), .B(OR4_514_Y), .C(OR4_205_Y), .D(
        OR4_68_Y), .Y(OR4_722_Y));
    OR4 OR4_172 (.A(sel_R_DATA_TEMPR32[10] ), .B(sel_R_DATA_TEMPR33[10] ), 
        .C(sel_R_DATA_TEMPR34[10] ), .D(sel_R_DATA_TEMPR35[10] ), .Y(
        OR4_172_Y));
    OR4 OR4_745 (.A(\SB_CORRECT[96] ), .B(\SB_CORRECT[97] ), .C(
        \SB_CORRECT[98] ), .D(\SB_CORRECT[99] ), .Y(OR4_745_Y));
    OR4 OR4_647 (.A(sel_R_DATA_TEMPR116[6] ), .B(sel_R_DATA_TEMPR117[6] ), 
        .C(sel_R_DATA_TEMPR118[6] ), .D(sel_R_DATA_TEMPR119[6] ), .Y(
        OR4_647_Y));
    OR4 OR4_1386 (.A(sel_R_DATA_TEMPR24[7] ), .B(sel_R_DATA_TEMPR25[7] ), .C(sel_R_DATA_TEMPR26[7] ), .D(sel_R_DATA_TEMPR27[7] ), .Y(OR4_1386_Y));
    OR4 OR4_975 (.A(sel_R_DATA_TEMPR64[0] ), .B(sel_R_DATA_TEMPR65[0] ), .C(sel_R_DATA_TEMPR66[0] ), .D(sel_R_DATA_TEMPR67[0] ), .Y(OR4_975_Y));
    OR4 OR4_1254 (.A(sel_R_DATA_TEMPR40[12] ), .B(sel_R_DATA_TEMPR41[12] ), 
        .C(sel_R_DATA_TEMPR42[12] ), .D(sel_R_DATA_TEMPR43[12] ), .Y(
        OR4_1254_Y));
    OR4 OR4_816 (.A(\SB_CORRECT[120] ), .B(\SB_CORRECT[121] ), 
        .C(\SB_CORRECT[122] ), .D(\SB_CORRECT[123] ), .Y(
        OR4_816_Y));
    AND4 \AND4SB_CORRECT[59]  (.A(sel_SB_CORRECT_NG[59] ), .B(
        \BLKY2_pipe[14] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[59] ));
    OR4 OR4_746 (.A(sel_R_DATA_TEMPR0[4] ), .B(sel_R_DATA_TEMPR1[4] ), .C(sel_R_DATA_TEMPR2[4] ), .D(sel_R_DATA_TEMPR3[4] ), .Y(OR4_746_Y));
    OR4 OR4_711 (.A(sel_R_DATA_TEMPR96[22] ), .B(sel_R_DATA_TEMPR97[22] ), 
        .C(sel_R_DATA_TEMPR98[22] ), .D(sel_R_DATA_TEMPR99[22] ), .Y(
        OR4_711_Y));
    OR4 OR4_585 (.A(\SB_CORRECT[108] ), .B(\SB_CORRECT[109] ), 
        .C(\SB_CORRECT[110] ), .D(\SB_CORRECT[111] ), .Y(
        OR4_585_Y));
    AND4 \AND4DB_DETECT[78]  (.A(sel_DB_DETECT_NG[78] ), .B(
        \BLKY2_pipe[19] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[78] ));
    OR4 OR4_926 (.A(sel_R_DATA_TEMPR44[29] ), .B(sel_R_DATA_TEMPR45[29] ), 
        .C(sel_R_DATA_TEMPR46[29] ), .D(sel_R_DATA_TEMPR47[29] ), .Y(
        OR4_926_Y));
    OR4 OR4_767 (.A(sel_R_DATA_TEMPR56[30] ), .B(sel_R_DATA_TEMPR57[30] ), 
        .C(sel_R_DATA_TEMPR58[30] ), .D(sel_R_DATA_TEMPR59[30] ), .Y(
        OR4_767_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%112%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R112C0 (.A_DOUT({
        nc408, nc409, nc410, nc411, nc412,int_R_DATA_TEMPR112[31] , 
       int_R_DATA_TEMPR112[30] ,int_R_DATA_TEMPR112[29] , 
       int_R_DATA_TEMPR112[28] ,int_R_DATA_TEMPR112[27] , 
       int_R_DATA_TEMPR112[26] ,int_R_DATA_TEMPR112[25] , 
       int_R_DATA_TEMPR112[24] ,int_R_DATA_TEMPR112[23] , 
       int_R_DATA_TEMPR112[22] ,int_R_DATA_TEMPR112[21] , 
       int_R_DATA_TEMPR112[20] ,int_R_DATA_TEMPR112[19] , 
       int_R_DATA_TEMPR112[18] ,int_R_DATA_TEMPR112[17] }), .B_DOUT({nc413, 
        nc414, nc415,int_R_DATA_TEMPR112[16] ,int_R_DATA_TEMPR112[15] , 
       int_R_DATA_TEMPR112[14] ,int_R_DATA_TEMPR112[13] , 
       int_R_DATA_TEMPR112[12] ,int_R_DATA_TEMPR112[11] , 
       int_R_DATA_TEMPR112[10] ,int_R_DATA_TEMPR112[9] , 
       int_R_DATA_TEMPR112[8] ,int_R_DATA_TEMPR112[7] , 
       int_R_DATA_TEMPR112[6] ,int_R_DATA_TEMPR112[5] , 
       int_R_DATA_TEMPR112[4] ,int_R_DATA_TEMPR112[3] , 
       int_R_DATA_TEMPR112[2] ,int_R_DATA_TEMPR112[1] , 
       int_R_DATA_TEMPR112[0] }), .DB_DETECT(int_DB_DETECT_NG[112] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[112] ), .ACCESS_BUSY(
        ACCESS_BUSY[112] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[28] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[28] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_255 (.A(sel_R_DATA_TEMPR124[18] ), .B(sel_R_DATA_TEMPR125[18] ), 
        .C(sel_R_DATA_TEMPR126[18] ), .D(sel_R_DATA_TEMPR127[18] ), .Y(
        OR4_255_Y));
    OR4 OR4_397 (.A(sel_R_DATA_TEMPR44[1] ), .B(sel_R_DATA_TEMPR45[1] ), .C(sel_R_DATA_TEMPR46[1] ), .D(sel_R_DATA_TEMPR47[1] ), .Y(OR4_397_Y));
    OR4 OR4_190 (.A(sel_R_DATA_TEMPR92[19] ), .B(sel_R_DATA_TEMPR93[19] ), 
        .C(sel_R_DATA_TEMPR94[19] ), .D(sel_R_DATA_TEMPR95[19] ), .Y(
        OR4_190_Y));
    OR4 OR4_1357 (.A(sel_R_DATA_TEMPR40[30] ), .B(sel_R_DATA_TEMPR41[30] ), 
        .C(sel_R_DATA_TEMPR42[30] ), .D(sel_R_DATA_TEMPR43[30] ), .Y(
        OR4_1357_Y));
    OR4 OR4_764 (.A(sel_R_DATA_TEMPR44[15] ), .B(sel_R_DATA_TEMPR45[15] ), 
        .C(sel_R_DATA_TEMPR46[15] ), .D(sel_R_DATA_TEMPR47[15] ), .Y(
        OR4_764_Y));
    OR4 OR4_625 (.A(sel_R_DATA_TEMPR64[21] ), .B(sel_R_DATA_TEMPR65[21] ), 
        .C(sel_R_DATA_TEMPR66[21] ), .D(sel_R_DATA_TEMPR67[21] ), .Y(
        OR4_625_Y));
    AND4 \AND4SB_CORRECT[17]  (.A(sel_SB_CORRECT_NG[17] ), .B(
        \BLKY2_pipe[4] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[17] ));
    OR4 OR4_852 (.A(OR4_1024_Y), .B(OR4_117_Y), .C(OR4_783_Y), .D(
        OR4_1007_Y), .Y(OR4_852_Y));
    OR4 OR4_538 (.A(sel_R_DATA_TEMPR36[19] ), .B(sel_R_DATA_TEMPR37[19] ), 
        .C(sel_R_DATA_TEMPR38[19] ), .D(sel_R_DATA_TEMPR39[19] ), .Y(
        OR4_538_Y));
    OR4 OR4_26 (.A(OR4_1230_Y), .B(OR4_96_Y), .C(OR4_1005_Y), .D(
        OR4_351_Y), .Y(OR4_26_Y));
    OR4 OR4_53 (.A(sel_R_DATA_TEMPR0[17] ), .B(sel_R_DATA_TEMPR1[17] ), .C(sel_R_DATA_TEMPR2[17] ), .D(sel_R_DATA_TEMPR3[17] ), .Y(OR4_53_Y));
    OR4 OR4_683 (.A(sel_R_DATA_TEMPR104[25] ), .B(sel_R_DATA_TEMPR105[25] ), 
        .C(sel_R_DATA_TEMPR106[25] ), .D(sel_R_DATA_TEMPR107[25] ), .Y(
        OR4_683_Y));
    AND4 \AND4SB_CORRECT[34]  (.A(sel_SB_CORRECT_NG[34] ), .B(
        \BLKY2_pipe[8] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[34] ));
    OR4 OR4_209 (.A(OR4_975_Y), .B(OR4_1213_Y), .C(OR4_1370_Y), .D(
        OR4_1167_Y), .Y(OR4_209_Y));
    OR4 OR4_798 (.A(\SB_CORRECT[100] ), .B(\SB_CORRECT[101] ), 
        .C(\SB_CORRECT[102] ), .D(\SB_CORRECT[103] ), .Y(
        OR4_798_Y));
    OR4 OR4_861 (.A(OR4_738_Y), .B(OR2_8_Y), .C(sel_R_DATA_TEMPR86[24] ), 
        .D(sel_R_DATA_TEMPR87[24] ), .Y(OR4_861_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%110%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R110C0 (.A_DOUT({
        nc416, nc417, nc418, nc419, nc420,int_R_DATA_TEMPR110[31] , 
       int_R_DATA_TEMPR110[30] ,int_R_DATA_TEMPR110[29] , 
       int_R_DATA_TEMPR110[28] ,int_R_DATA_TEMPR110[27] , 
       int_R_DATA_TEMPR110[26] ,int_R_DATA_TEMPR110[25] , 
       int_R_DATA_TEMPR110[24] ,int_R_DATA_TEMPR110[23] , 
       int_R_DATA_TEMPR110[22] ,int_R_DATA_TEMPR110[21] , 
       int_R_DATA_TEMPR110[20] ,int_R_DATA_TEMPR110[19] , 
       int_R_DATA_TEMPR110[18] ,int_R_DATA_TEMPR110[17] }), .B_DOUT({nc421, 
        nc422, nc423,int_R_DATA_TEMPR110[16] ,int_R_DATA_TEMPR110[15] , 
       int_R_DATA_TEMPR110[14] ,int_R_DATA_TEMPR110[13] , 
       int_R_DATA_TEMPR110[12] ,int_R_DATA_TEMPR110[11] , 
       int_R_DATA_TEMPR110[10] ,int_R_DATA_TEMPR110[9] , 
       int_R_DATA_TEMPR110[8] ,int_R_DATA_TEMPR110[7] , 
       int_R_DATA_TEMPR110[6] ,int_R_DATA_TEMPR110[5] , 
       int_R_DATA_TEMPR110[4] ,int_R_DATA_TEMPR110[3] , 
       int_R_DATA_TEMPR110[2] ,int_R_DATA_TEMPR110[1] , 
       int_R_DATA_TEMPR110[0] }), .DB_DETECT(int_DB_DETECT_NG[110] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[110] ), .ACCESS_BUSY(
        ACCESS_BUSY[110] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[27] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[27] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%113%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R113C0 (.A_DOUT({
        nc424, nc425, nc426, nc427, nc428,int_R_DATA_TEMPR113[31] , 
       int_R_DATA_TEMPR113[30] ,int_R_DATA_TEMPR113[29] , 
       int_R_DATA_TEMPR113[28] ,int_R_DATA_TEMPR113[27] , 
       int_R_DATA_TEMPR113[26] ,int_R_DATA_TEMPR113[25] , 
       int_R_DATA_TEMPR113[24] ,int_R_DATA_TEMPR113[23] , 
       int_R_DATA_TEMPR113[22] ,int_R_DATA_TEMPR113[21] , 
       int_R_DATA_TEMPR113[20] ,int_R_DATA_TEMPR113[19] , 
       int_R_DATA_TEMPR113[18] ,int_R_DATA_TEMPR113[17] }), .B_DOUT({nc429, 
        nc430, nc431,int_R_DATA_TEMPR113[16] ,int_R_DATA_TEMPR113[15] , 
       int_R_DATA_TEMPR113[14] ,int_R_DATA_TEMPR113[13] , 
       int_R_DATA_TEMPR113[12] ,int_R_DATA_TEMPR113[11] , 
       int_R_DATA_TEMPR113[10] ,int_R_DATA_TEMPR113[9] , 
       int_R_DATA_TEMPR113[8] ,int_R_DATA_TEMPR113[7] , 
       int_R_DATA_TEMPR113[6] ,int_R_DATA_TEMPR113[5] , 
       int_R_DATA_TEMPR113[4] ,int_R_DATA_TEMPR113[3] , 
       int_R_DATA_TEMPR113[2] ,int_R_DATA_TEMPR113[1] , 
       int_R_DATA_TEMPR113[0] }), .DB_DETECT(int_DB_DETECT_NG[113] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[113] ), .ACCESS_BUSY(
        ACCESS_BUSY[113] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[28] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[28] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_516 (.A(sel_R_DATA_TEMPR116[9] ), .B(sel_R_DATA_TEMPR117[9] ), 
        .C(sel_R_DATA_TEMPR118[9] ), .D(sel_R_DATA_TEMPR119[9] ), .Y(
        OR4_516_Y));
    AND4 \AND4SB_CORRECT[3]  (.A(sel_SB_CORRECT_NG[3] ), .B(
        \BLKY2_pipe[0] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[3] ));
    OR4 OR4_279 (.A(sel_R_DATA_TEMPR108[15] ), .B(sel_R_DATA_TEMPR109[15] ), 
        .C(sel_R_DATA_TEMPR110[15] ), .D(sel_R_DATA_TEMPR111[15] ), .Y(
        OR4_279_Y));
    OR4 OR4_1267 (.A(sel_R_DATA_TEMPR48[2] ), .B(sel_R_DATA_TEMPR49[2] ), .C(sel_R_DATA_TEMPR50[2] ), .D(sel_R_DATA_TEMPR51[2] ), .Y(OR4_1267_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[30]  (.D(\BLKY2[30] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[30] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%83%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R83C0 (.A_DOUT({
        nc432, nc433, nc434, nc435, nc436,int_R_DATA_TEMPR83[31] , 
       int_R_DATA_TEMPR83[30] ,int_R_DATA_TEMPR83[29] , 
       int_R_DATA_TEMPR83[28] ,int_R_DATA_TEMPR83[27] , 
       int_R_DATA_TEMPR83[26] ,int_R_DATA_TEMPR83[25] , 
       int_R_DATA_TEMPR83[24] ,int_R_DATA_TEMPR83[23] , 
       int_R_DATA_TEMPR83[22] ,int_R_DATA_TEMPR83[21] , 
       int_R_DATA_TEMPR83[20] ,int_R_DATA_TEMPR83[19] , 
       int_R_DATA_TEMPR83[18] ,int_R_DATA_TEMPR83[17] }), .B_DOUT({nc437, 
        nc438, nc439,int_R_DATA_TEMPR83[16] ,int_R_DATA_TEMPR83[15] , 
       int_R_DATA_TEMPR83[14] ,int_R_DATA_TEMPR83[13] , 
       int_R_DATA_TEMPR83[12] ,int_R_DATA_TEMPR83[11] , 
       int_R_DATA_TEMPR83[10] ,int_R_DATA_TEMPR83[9] ,int_R_DATA_TEMPR83[8] , 
       int_R_DATA_TEMPR83[7] ,int_R_DATA_TEMPR83[6] ,int_R_DATA_TEMPR83[5] , 
       int_R_DATA_TEMPR83[4] ,int_R_DATA_TEMPR83[3] ,int_R_DATA_TEMPR83[2] , 
       int_R_DATA_TEMPR83[1] ,int_R_DATA_TEMPR83[0] }), .DB_DETECT( int_DB_DETECT_NG[83] ), .SB_CORRECT(int_SB_CORRECT_NG[83] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[83] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[20] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[20] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_436 (.A(OR4_726_Y), .B(OR4_1237_Y), .C(OR4_507_Y), .D(
        OR4_719_Y), .Y(OR4_436_Y));
    OR4 OR4_453 (.A(OR4_1372_Y), .B(OR4_238_Y), .C(OR4_1160_Y), .D(
        OR4_501_Y), .Y(OR4_453_Y));
    OR4 OR4_89 (.A(sel_R_DATA_TEMPR8[11] ), .B(sel_R_DATA_TEMPR9[11] ), .C(sel_R_DATA_TEMPR10[11] ), .D(sel_R_DATA_TEMPR11[11] ), .Y(OR4_89_Y));
    OR4 OR4_1104 (.A(sel_R_DATA_TEMPR24[17] ), .B(sel_R_DATA_TEMPR25[17] ), 
        .C(sel_R_DATA_TEMPR26[17] ), .D(sel_R_DATA_TEMPR27[17] ), .Y(
        OR4_1104_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%91%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R91C0 (.A_DOUT({
        nc440, nc441, nc442, nc443, nc444,int_R_DATA_TEMPR91[31] , 
       int_R_DATA_TEMPR91[30] ,int_R_DATA_TEMPR91[29] , 
       int_R_DATA_TEMPR91[28] ,int_R_DATA_TEMPR91[27] , 
       int_R_DATA_TEMPR91[26] ,int_R_DATA_TEMPR91[25] , 
       int_R_DATA_TEMPR91[24] ,int_R_DATA_TEMPR91[23] , 
       int_R_DATA_TEMPR91[22] ,int_R_DATA_TEMPR91[21] , 
       int_R_DATA_TEMPR91[20] ,int_R_DATA_TEMPR91[19] , 
       int_R_DATA_TEMPR91[18] ,int_R_DATA_TEMPR91[17] }), .B_DOUT({nc445, 
        nc446, nc447,int_R_DATA_TEMPR91[16] ,int_R_DATA_TEMPR91[15] , 
       int_R_DATA_TEMPR91[14] ,int_R_DATA_TEMPR91[13] , 
       int_R_DATA_TEMPR91[12] ,int_R_DATA_TEMPR91[11] , 
       int_R_DATA_TEMPR91[10] ,int_R_DATA_TEMPR91[9] ,int_R_DATA_TEMPR91[8] , 
       int_R_DATA_TEMPR91[7] ,int_R_DATA_TEMPR91[6] ,int_R_DATA_TEMPR91[5] , 
       int_R_DATA_TEMPR91[4] ,int_R_DATA_TEMPR91[3] ,int_R_DATA_TEMPR91[2] , 
       int_R_DATA_TEMPR91[1] ,int_R_DATA_TEMPR91[0] }), .DB_DETECT( int_DB_DETECT_NG[91] ), .SB_CORRECT(int_SB_CORRECT_NG[91] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[91] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[22] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[22] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_897 (.A(sel_R_DATA_TEMPR40[13] ), .B(sel_R_DATA_TEMPR41[13] ), 
        .C(sel_R_DATA_TEMPR42[13] ), .D(sel_R_DATA_TEMPR43[13] ), .Y(
        OR4_897_Y));
    OR4 OR4_651 (.A(sel_R_DATA_TEMPR76[10] ), .B(sel_R_DATA_TEMPR77[10] ), 
        .C(sel_R_DATA_TEMPR78[10] ), .D(sel_R_DATA_TEMPR79[10] ), .Y(
        OR4_651_Y));
    OR4 OR4_198 (.A(sel_R_DATA_TEMPR28[28] ), .B(sel_R_DATA_TEMPR29[28] ), 
        .C(sel_R_DATA_TEMPR30[28] ), .D(sel_R_DATA_TEMPR31[28] ), .Y(
        OR4_198_Y));
    OR4 OR4_1078 (.A(\DB_DETECT[0] ), .B(\DB_DETECT[1] ), .C(
        \DB_DETECT[2] ), .D(\DB_DETECT[3] ), .Y(OR4_1078_Y));
    OR4 OR4_994 (.A(\SB_CORRECT[112] ), .B(\SB_CORRECT[113] ), 
        .C(\SB_CORRECT[114] ), .D(\SB_CORRECT[115] ), .Y(
        OR4_994_Y));
    OR4 OR4_989 (.A(sel_R_DATA_TEMPR40[8] ), .B(sel_R_DATA_TEMPR41[8] ), .C(sel_R_DATA_TEMPR42[8] ), .D(sel_R_DATA_TEMPR43[8] ), .Y(OR4_989_Y));
    OR4 OR4_980 (.A(sel_R_DATA_TEMPR112[13] ), .B(sel_R_DATA_TEMPR113[13] ), 
        .C(sel_R_DATA_TEMPR114[13] ), .D(sel_R_DATA_TEMPR115[13] ), .Y(
        OR4_980_Y));
    OR4 OR4_809 (.A(sel_R_DATA_TEMPR116[30] ), .B(sel_R_DATA_TEMPR117[30] ), 
        .C(sel_R_DATA_TEMPR118[30] ), .D(sel_R_DATA_TEMPR119[30] ), .Y(
        OR4_809_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[3]  (.A(CFG3_5_Y), .B(CFG3_12_Y)
        , .Y(\BLKX2[3] ));
    OR4 OR4_258 (.A(sel_R_DATA_TEMPR76[28] ), .B(sel_R_DATA_TEMPR77[28] ), 
        .C(sel_R_DATA_TEMPR78[28] ), .D(sel_R_DATA_TEMPR79[28] ), .Y(
        OR4_258_Y));
    OR4 OR4_1364 (.A(sel_R_DATA_TEMPR16[25] ), .B(sel_R_DATA_TEMPR17[25] ), 
        .C(sel_R_DATA_TEMPR18[25] ), .D(sel_R_DATA_TEMPR19[25] ), .Y(
        OR4_1364_Y));
    OR4 \OR4_R_DATA[21]  (.A(OR4_1279_Y), .B(OR4_1217_Y), .C(
        OR4_1244_Y), .D(OR4_785_Y), .Y(R_DATA[21]));
    OR4 OR4_1123 (.A(sel_R_DATA_TEMPR88[16] ), .B(sel_R_DATA_TEMPR89[16] ), 
        .C(sel_R_DATA_TEMPR90[16] ), .D(sel_R_DATA_TEMPR91[16] ), .Y(
        OR4_1123_Y));
    AND4 \AND4SB_CORRECT[106]  (.A(sel_SB_CORRECT_NG[106] ), .B(
        \BLKY2_pipe[26] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[106] ));
    OR4 OR4_620 (.A(sel_R_DATA_TEMPR64[8] ), .B(sel_R_DATA_TEMPR65[8] ), .C(sel_R_DATA_TEMPR66[8] ), .D(sel_R_DATA_TEMPR67[8] ), .Y(OR4_620_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[27]  (.A(CFG3_5_Y), .B(CFG3_7_Y)
        , .Y(\BLKX2[27] ));
    OR4 OR4_1345 (.A(OR4_1182_Y), .B(OR4_52_Y), .C(OR4_958_Y), .D(
        OR4_311_Y), .Y(OR4_1345_Y));
    OR4 OR4_879 (.A(\DB_DETECT[124] ), .B(\DB_DETECT[125] ), .C(
        \DB_DETECT[126] ), .D(\DB_DETECT[127] ), .Y(OR4_879_Y));
    OR4 OR4_183 (.A(sel_R_DATA_TEMPR44[13] ), .B(sel_R_DATA_TEMPR45[13] ), 
        .C(sel_R_DATA_TEMPR46[13] ), .D(sel_R_DATA_TEMPR47[13] ), .Y(
        OR4_183_Y));
    OR4 OR4_1111 (.A(OR4_1367_Y), .B(OR4_465_Y), .C(OR4_1126_Y), .D(
        OR4_1358_Y), .Y(OR4_1111_Y));
    AND4 \AND4SB_CORRECT[103]  (.A(sel_SB_CORRECT_NG[103] ), .B(
        \BLKY2_pipe[25] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[103] ));
    OR4 OR4_332 (.A(sel_R_DATA_TEMPR72[24] ), .B(sel_R_DATA_TEMPR73[24] ), 
        .C(sel_R_DATA_TEMPR74[24] ), .D(sel_R_DATA_TEMPR75[24] ), .Y(
        OR4_332_Y));
    AND4 \AND4DB_DETECT[40]  (.A(sel_DB_DETECT_NG[40] ), .B(
        \BLKY2_pipe[10] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[40] ));
    AND4 \AND4DB_DETECT[9]  (.A(sel_DB_DETECT_NG[9] ), .B(
        \BLKY2_pipe[2] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[9] ));
    OR4 OR4_13 (.A(sel_R_DATA_TEMPR16[0] ), .B(sel_R_DATA_TEMPR17[0] ), .C(sel_R_DATA_TEMPR18[0] ), .D(sel_R_DATA_TEMPR19[0] ), .Y(OR4_13_Y));
    OR4 OR4_247 (.A(sel_R_DATA_TEMPR32[19] ), .B(sel_R_DATA_TEMPR33[19] ), 
        .C(sel_R_DATA_TEMPR34[19] ), .D(sel_R_DATA_TEMPR35[19] ), .Y(
        OR4_247_Y));
    OR4 OR4_1208 (.A(OR4_30_Y), .B(OR4_892_Y), .C(OR4_1115_Y), .D(
        OR4_217_Y), .Y(OR4_1208_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_3 (.A(R_EN), .B(R_ADDR[15]), .C(
        R_ADDR[14]), .Y(CFG3_3_Y));
    OR4 OR4_518 (.A(OR4_1361_Y), .B(OR4_865_Y), .C(OR4_59_Y), .D(
        OR4_650_Y), .Y(OR4_518_Y));
    OR4 OR4_147 (.A(sel_R_DATA_TEMPR96[11] ), .B(sel_R_DATA_TEMPR97[11] ), 
        .C(sel_R_DATA_TEMPR98[11] ), .D(sel_R_DATA_TEMPR99[11] ), .Y(
        OR4_147_Y));
    OR4 OR4_327 (.A(sel_R_DATA_TEMPR36[22] ), .B(sel_R_DATA_TEMPR37[22] ), 
        .C(sel_R_DATA_TEMPR38[22] ), .D(sel_R_DATA_TEMPR39[22] ), .Y(
        OR4_327_Y));
    OR4 OR4_120 (.A(sel_R_DATA_TEMPR104[26] ), .B(sel_R_DATA_TEMPR105[26] ), 
        .C(sel_R_DATA_TEMPR106[26] ), .D(sel_R_DATA_TEMPR107[26] ), .Y(
        OR4_120_Y));
    INV \INVBLKY1[0]  (.A(R_ADDR[10]), .Y(\BLKY1[0] ));
    OR4 OR4_51 (.A(OR4_617_Y), .B(OR4_872_Y), .C(OR4_423_Y), .D(
        OR4_1145_Y), .Y(OR4_51_Y));
    OR4 OR4_967 (.A(sel_R_DATA_TEMPR0[27] ), .B(sel_R_DATA_TEMPR1[27] ), .C(sel_R_DATA_TEMPR2[27] ), .D(sel_R_DATA_TEMPR3[27] ), .Y(OR4_967_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[10]  (.D(\BLKY2[10] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[10] ));
    DFN1E1 \DFN1E1BLKY2_pipe[26]  (.D(\BLKY2[26] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[26] ));
    OR2 OR2_2 (.A(sel_R_DATA_TEMPR84[25] ), .B(sel_R_DATA_TEMPR85[25] ), .Y(
        OR2_2_Y));
    AND4 \AND4DB_DETECT[8]  (.A(sel_DB_DETECT_NG[8] ), .B(
        \BLKY2_pipe[2] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[8] ));
    OR4 \OR4_R_DATA[20]  (.A(OR4_1010_Y), .B(OR4_1338_Y), .C(OR4_567_Y)
        , .D(OR4_44_Y), .Y(R_DATA[20]));
    OR4 OR4_1184 (.A(\DB_DETECT[112] ), .B(\DB_DETECT[113] ), .C(
        \DB_DETECT[114] ), .D(\DB_DETECT[115] ), .Y(OR4_1184_Y));
    AND4 \AND4DB_DETECT[93]  (.A(sel_DB_DETECT_NG[93] ), .B(
        \BLKY2_pipe[23] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[93] ));
    OR4 OR4_1236 (.A(sel_R_DATA_TEMPR104[30] ), .B(sel_R_DATA_TEMPR105[30] ), 
        .C(sel_R_DATA_TEMPR106[30] ), .D(sel_R_DATA_TEMPR107[30] ), .Y(
        OR4_1236_Y));
    OR4 OR4_728 (.A(sel_R_DATA_TEMPR40[16] ), .B(sel_R_DATA_TEMPR41[16] ), 
        .C(sel_R_DATA_TEMPR42[16] ), .D(sel_R_DATA_TEMPR43[16] ), .Y(
        OR4_728_Y));
    OR4 OR4_707 (.A(sel_R_DATA_TEMPR64[29] ), .B(sel_R_DATA_TEMPR65[29] ), 
        .C(sel_R_DATA_TEMPR66[29] ), .D(sel_R_DATA_TEMPR67[29] ), .Y(
        OR4_707_Y));
    OR4 OR4_1297 (.A(sel_R_DATA_TEMPR88[7] ), .B(sel_R_DATA_TEMPR89[7] ), .C(sel_R_DATA_TEMPR90[7] ), .D(sel_R_DATA_TEMPR91[7] ), .Y(OR4_1297_Y));
    OR4 OR4_704 (.A(sel_R_DATA_TEMPR92[25] ), .B(sel_R_DATA_TEMPR93[25] ), 
        .C(sel_R_DATA_TEMPR94[25] ), .D(sel_R_DATA_TEMPR95[25] ), .Y(
        OR4_704_Y));
    OR4 OR4_1369 (.A(sel_R_DATA_TEMPR64[20] ), .B(sel_R_DATA_TEMPR65[20] ), 
        .C(sel_R_DATA_TEMPR66[20] ), .D(sel_R_DATA_TEMPR67[20] ), .Y(
        OR4_1369_Y));
    OR4 OR4_20 (.A(sel_R_DATA_TEMPR100[25] ), .B(sel_R_DATA_TEMPR101[25] ), 
        .C(sel_R_DATA_TEMPR102[25] ), .D(sel_R_DATA_TEMPR103[25] ), .Y(
        OR4_20_Y));
    OR4 OR4_1338 (.A(OR4_150_Y), .B(OR4_687_Y), .C(OR4_1154_Y), .D(
        OR4_633_Y), .Y(OR4_1338_Y));
    OR4 OR4_743 (.A(sel_R_DATA_TEMPR100[9] ), .B(sel_R_DATA_TEMPR101[9] ), 
        .C(sel_R_DATA_TEMPR102[9] ), .D(sel_R_DATA_TEMPR103[9] ), .Y(
        OR4_743_Y));
    OR4 OR4_1060 (.A(sel_R_DATA_TEMPR64[2] ), .B(sel_R_DATA_TEMPR65[2] ), .C(sel_R_DATA_TEMPR66[2] ), .D(sel_R_DATA_TEMPR67[2] ), .Y(OR4_1060_Y));
    OR4 OR4_777 (.A(sel_R_DATA_TEMPR4[0] ), .B(sel_R_DATA_TEMPR5[0] ), .C(sel_R_DATA_TEMPR6[0] ), .D(sel_R_DATA_TEMPR7[0] ), .Y(OR4_777_Y));
    AND4 \AND4DB_DETECT[63]  (.A(sel_DB_DETECT_NG[63] ), .B(
        \BLKY2_pipe[15] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[63] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%4%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R4C0 (.A_DOUT({
        nc448, nc449, nc450, nc451, nc452,int_R_DATA_TEMPR4[31] , 
       int_R_DATA_TEMPR4[30] ,int_R_DATA_TEMPR4[29] ,int_R_DATA_TEMPR4[28] , 
       int_R_DATA_TEMPR4[27] ,int_R_DATA_TEMPR4[26] ,int_R_DATA_TEMPR4[25] , 
       int_R_DATA_TEMPR4[24] ,int_R_DATA_TEMPR4[23] ,int_R_DATA_TEMPR4[22] , 
       int_R_DATA_TEMPR4[21] ,int_R_DATA_TEMPR4[20] ,int_R_DATA_TEMPR4[19] , 
       int_R_DATA_TEMPR4[18] ,int_R_DATA_TEMPR4[17] }), .B_DOUT({nc453, 
        nc454, nc455,int_R_DATA_TEMPR4[16] ,int_R_DATA_TEMPR4[15] , 
       int_R_DATA_TEMPR4[14] ,int_R_DATA_TEMPR4[13] ,int_R_DATA_TEMPR4[12] , 
       int_R_DATA_TEMPR4[11] ,int_R_DATA_TEMPR4[10] ,int_R_DATA_TEMPR4[9] , 
       int_R_DATA_TEMPR4[8] ,int_R_DATA_TEMPR4[7] ,int_R_DATA_TEMPR4[6] , 
       int_R_DATA_TEMPR4[5] ,int_R_DATA_TEMPR4[4] ,int_R_DATA_TEMPR4[3] , 
       int_R_DATA_TEMPR4[2] ,int_R_DATA_TEMPR4[1] ,int_R_DATA_TEMPR4[0] }), 
        .DB_DETECT(int_DB_DETECT_NG[4] ), .SB_CORRECT( int_SB_CORRECT_NG[4] ), .ACCESS_BUSY(\ACCESS_BUSY[4] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[1] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_416 (.A(sel_R_DATA_TEMPR32[0] ), .B(sel_R_DATA_TEMPR33[0] ), .C(sel_R_DATA_TEMPR34[0] ), .D(sel_R_DATA_TEMPR35[0] ), .Y(OR4_416_Y));
    OR4 \OR4_R_DATA[26]  (.A(OR4_525_Y), .B(OR4_1286_Y), .C(OR4_134_Y), 
        .D(OR4_216_Y), .Y(R_DATA[26]));
    OR4 OR4_774 (.A(sel_R_DATA_TEMPR100[5] ), .B(sel_R_DATA_TEMPR101[5] ), 
        .C(sel_R_DATA_TEMPR102[5] ), .D(sel_R_DATA_TEMPR103[5] ), .Y(
        OR4_774_Y));
    AND4 \AND4SB_CORRECT[22]  (.A(sel_SB_CORRECT_NG[22] ), .B(
        \BLKY2_pipe[5] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[22] ));
    OR4 OR4_244 (.A(sel_R_DATA_TEMPR80[5] ), .B(sel_R_DATA_TEMPR81[5] ), .C(sel_R_DATA_TEMPR82[5] ), .D(sel_R_DATA_TEMPR83[5] ), .Y(OR4_244_Y));
    OR4 OR4_1356 (.A(sel_R_DATA_TEMPR32[8] ), .B(sel_R_DATA_TEMPR33[8] ), .C(sel_R_DATA_TEMPR34[8] ), .D(sel_R_DATA_TEMPR35[8] ), .Y(OR4_1356_Y));
    OR4 OR4_801 (.A(sel_R_DATA_TEMPR16[3] ), .B(sel_R_DATA_TEMPR17[3] ), .C(sel_R_DATA_TEMPR18[3] ), .D(sel_R_DATA_TEMPR19[3] ), .Y(OR4_801_Y));
    AND4 \AND4DB_DETECT[79]  (.A(sel_DB_DETECT_NG[79] ), .B(
        \BLKY2_pipe[19] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[79] ));
    OR4 OR4_1288 (.A(sel_R_DATA_TEMPR20[14] ), .B(sel_R_DATA_TEMPR21[14] ), 
        .C(sel_R_DATA_TEMPR22[14] ), .D(sel_R_DATA_TEMPR23[14] ), .Y(
        OR4_1288_Y));
    OR4 OR4_27 (.A(sel_R_DATA_TEMPR20[12] ), .B(sel_R_DATA_TEMPR21[12] ), .C(sel_R_DATA_TEMPR22[12] ), .D(sel_R_DATA_TEMPR23[12] ), .Y(OR4_27_Y));
    AND4 \AND4SB_CORRECT[78]  (.A(sel_SB_CORRECT_NG[78] ), .B(
        \BLKY2_pipe[19] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[78] ));
    OR4 OR4_82 (.A(sel_R_DATA_TEMPR104[13] ), .B(sel_R_DATA_TEMPR105[13] ), 
        .C(sel_R_DATA_TEMPR106[13] ), .D(sel_R_DATA_TEMPR107[13] ), .Y(
        OR4_82_Y));
    OR4 OR4_827 (.A(sel_R_DATA_TEMPR108[20] ), .B(sel_R_DATA_TEMPR109[20] ), 
        .C(sel_R_DATA_TEMPR110[20] ), .D(sel_R_DATA_TEMPR111[20] ), .Y(
        OR4_827_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%44%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R44C0 (.A_DOUT({
        nc456, nc457, nc458, nc459, nc460,int_R_DATA_TEMPR44[31] , 
       int_R_DATA_TEMPR44[30] ,int_R_DATA_TEMPR44[29] , 
       int_R_DATA_TEMPR44[28] ,int_R_DATA_TEMPR44[27] , 
       int_R_DATA_TEMPR44[26] ,int_R_DATA_TEMPR44[25] , 
       int_R_DATA_TEMPR44[24] ,int_R_DATA_TEMPR44[23] , 
       int_R_DATA_TEMPR44[22] ,int_R_DATA_TEMPR44[21] , 
       int_R_DATA_TEMPR44[20] ,int_R_DATA_TEMPR44[19] , 
       int_R_DATA_TEMPR44[18] ,int_R_DATA_TEMPR44[17] }), .B_DOUT({nc461, 
        nc462, nc463,int_R_DATA_TEMPR44[16] ,int_R_DATA_TEMPR44[15] , 
       int_R_DATA_TEMPR44[14] ,int_R_DATA_TEMPR44[13] , 
       int_R_DATA_TEMPR44[12] ,int_R_DATA_TEMPR44[11] , 
       int_R_DATA_TEMPR44[10] ,int_R_DATA_TEMPR44[9] ,int_R_DATA_TEMPR44[8] , 
       int_R_DATA_TEMPR44[7] ,int_R_DATA_TEMPR44[6] ,int_R_DATA_TEMPR44[5] , 
       int_R_DATA_TEMPR44[4] ,int_R_DATA_TEMPR44[3] ,int_R_DATA_TEMPR44[2] , 
       int_R_DATA_TEMPR44[1] ,int_R_DATA_TEMPR44[0] }), .DB_DETECT( int_DB_DETECT_NG[44] ), .SB_CORRECT(int_SB_CORRECT_NG[44] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[44] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[11] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[11] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_128 (.A(sel_R_DATA_TEMPR100[28] ), .B(sel_R_DATA_TEMPR101[28] ), 
        .C(sel_R_DATA_TEMPR102[28] ), .D(sel_R_DATA_TEMPR103[28] ), .Y(
        OR4_128_Y));
    OR4 OR4_230 (.A(sel_R_DATA_TEMPR104[12] ), .B(sel_R_DATA_TEMPR105[12] ), 
        .C(sel_R_DATA_TEMPR106[12] ), .D(sel_R_DATA_TEMPR107[12] ), .Y(
        OR4_230_Y));
    OR4 OR4_924 (.A(sel_R_DATA_TEMPR64[26] ), .B(sel_R_DATA_TEMPR65[26] ), 
        .C(sel_R_DATA_TEMPR66[26] ), .D(sel_R_DATA_TEMPR67[26] ), .Y(
        OR4_924_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%105%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R105C0 (.A_DOUT({
        nc464, nc465, nc466, nc467, nc468,int_R_DATA_TEMPR105[31] , 
       int_R_DATA_TEMPR105[30] ,int_R_DATA_TEMPR105[29] , 
       int_R_DATA_TEMPR105[28] ,int_R_DATA_TEMPR105[27] , 
       int_R_DATA_TEMPR105[26] ,int_R_DATA_TEMPR105[25] , 
       int_R_DATA_TEMPR105[24] ,int_R_DATA_TEMPR105[23] , 
       int_R_DATA_TEMPR105[22] ,int_R_DATA_TEMPR105[21] , 
       int_R_DATA_TEMPR105[20] ,int_R_DATA_TEMPR105[19] , 
       int_R_DATA_TEMPR105[18] ,int_R_DATA_TEMPR105[17] }), .B_DOUT({nc469, 
        nc470, nc471,int_R_DATA_TEMPR105[16] ,int_R_DATA_TEMPR105[15] , 
       int_R_DATA_TEMPR105[14] ,int_R_DATA_TEMPR105[13] , 
       int_R_DATA_TEMPR105[12] ,int_R_DATA_TEMPR105[11] , 
       int_R_DATA_TEMPR105[10] ,int_R_DATA_TEMPR105[9] , 
       int_R_DATA_TEMPR105[8] ,int_R_DATA_TEMPR105[7] , 
       int_R_DATA_TEMPR105[6] ,int_R_DATA_TEMPR105[5] , 
       int_R_DATA_TEMPR105[4] ,int_R_DATA_TEMPR105[3] , 
       int_R_DATA_TEMPR105[2] ,int_R_DATA_TEMPR105[1] , 
       int_R_DATA_TEMPR105[0] }), .DB_DETECT(int_DB_DETECT_NG[105] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[105] ), .ACCESS_BUSY(
        ACCESS_BUSY[105] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[26] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[26] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1015 (.A(sel_R_DATA_TEMPR88[22] ), .B(sel_R_DATA_TEMPR89[22] ), 
        .C(sel_R_DATA_TEMPR90[22] ), .D(sel_R_DATA_TEMPR91[22] ), .Y(
        OR4_1015_Y));
    OR4 OR4_537 (.A(sel_R_DATA_TEMPR72[13] ), .B(sel_R_DATA_TEMPR73[13] ), 
        .C(sel_R_DATA_TEMPR74[13] ), .D(sel_R_DATA_TEMPR75[13] ), .Y(
        OR4_537_Y));
    OR4 OR4_880 (.A(\SB_CORRECT[116] ), .B(\SB_CORRECT[117] ), 
        .C(\SB_CORRECT[118] ), .D(\SB_CORRECT[119] ), .Y(
        OR4_880_Y));
    OR4 OR4_871 (.A(sel_R_DATA_TEMPR124[8] ), .B(sel_R_DATA_TEMPR125[8] ), 
        .C(sel_R_DATA_TEMPR126[8] ), .D(sel_R_DATA_TEMPR127[8] ), .Y(
        OR4_871_Y));
    OR4 OR4_182 (.A(sel_R_DATA_TEMPR80[31] ), .B(sel_R_DATA_TEMPR81[31] ), 
        .C(sel_R_DATA_TEMPR82[31] ), .D(sel_R_DATA_TEMPR83[31] ), .Y(
        OR4_182_Y));
    OR4 OR4_465 (.A(sel_R_DATA_TEMPR52[26] ), .B(sel_R_DATA_TEMPR53[26] ), 
        .C(sel_R_DATA_TEMPR54[26] ), .D(sel_R_DATA_TEMPR55[26] ), .Y(
        OR4_465_Y));
    OR4 OR4_312 (.A(sel_R_DATA_TEMPR88[27] ), .B(sel_R_DATA_TEMPR89[27] ), 
        .C(sel_R_DATA_TEMPR90[27] ), .D(sel_R_DATA_TEMPR91[27] ), .Y(
        OR4_312_Y));
    OR4 OR4_551 (.A(sel_R_DATA_TEMPR24[9] ), .B(sel_R_DATA_TEMPR25[9] ), .C(sel_R_DATA_TEMPR26[9] ), .D(sel_R_DATA_TEMPR27[9] ), .Y(OR4_551_Y));
    OR4 OR4_64 (.A(OR4_274_Y), .B(OR4_252_Y), .C(OR4_224_Y), .D(
        OR4_876_Y), .Y(OR4_64_Y));
    OR4 OR4_1105 (.A(sel_R_DATA_TEMPR80[15] ), .B(sel_R_DATA_TEMPR81[15] ), 
        .C(sel_R_DATA_TEMPR82[15] ), .D(sel_R_DATA_TEMPR83[15] ), .Y(
        OR4_1105_Y));
    OR4 OR4_1077 (.A(sel_R_DATA_TEMPR16[6] ), .B(sel_R_DATA_TEMPR17[6] ), .C(sel_R_DATA_TEMPR18[6] ), .D(sel_R_DATA_TEMPR19[6] ), .Y(OR4_1077_Y));
    OR4 OR4_985 (.A(sel_R_DATA_TEMPR64[5] ), .B(sel_R_DATA_TEMPR65[5] ), .C(sel_R_DATA_TEMPR66[5] ), .D(sel_R_DATA_TEMPR67[5] ), .Y(OR4_985_Y));
    OR4 OR4_11 (.A(sel_R_DATA_TEMPR28[16] ), .B(sel_R_DATA_TEMPR29[16] ), .C(sel_R_DATA_TEMPR30[16] ), .D(sel_R_DATA_TEMPR31[16] ), .Y(OR4_11_Y));
    OR4 OR4_1039 (.A(sel_R_DATA_TEMPR56[13] ), .B(sel_R_DATA_TEMPR57[13] ), 
        .C(sel_R_DATA_TEMPR58[13] ), .D(sel_R_DATA_TEMPR59[13] ), .Y(
        OR4_1039_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%18%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R18C0 (.A_DOUT({
        nc472, nc473, nc474, nc475, nc476,int_R_DATA_TEMPR18[31] , 
       int_R_DATA_TEMPR18[30] ,int_R_DATA_TEMPR18[29] , 
       int_R_DATA_TEMPR18[28] ,int_R_DATA_TEMPR18[27] , 
       int_R_DATA_TEMPR18[26] ,int_R_DATA_TEMPR18[25] , 
       int_R_DATA_TEMPR18[24] ,int_R_DATA_TEMPR18[23] , 
       int_R_DATA_TEMPR18[22] ,int_R_DATA_TEMPR18[21] , 
       int_R_DATA_TEMPR18[20] ,int_R_DATA_TEMPR18[19] , 
       int_R_DATA_TEMPR18[18] ,int_R_DATA_TEMPR18[17] }), .B_DOUT({nc477, 
        nc478, nc479,int_R_DATA_TEMPR18[16] ,int_R_DATA_TEMPR18[15] , 
       int_R_DATA_TEMPR18[14] ,int_R_DATA_TEMPR18[13] , 
       int_R_DATA_TEMPR18[12] ,int_R_DATA_TEMPR18[11] , 
       int_R_DATA_TEMPR18[10] ,int_R_DATA_TEMPR18[9] ,int_R_DATA_TEMPR18[8] , 
       int_R_DATA_TEMPR18[7] ,int_R_DATA_TEMPR18[6] ,int_R_DATA_TEMPR18[5] , 
       int_R_DATA_TEMPR18[4] ,int_R_DATA_TEMPR18[3] ,int_R_DATA_TEMPR18[2] , 
       int_R_DATA_TEMPR18[1] ,int_R_DATA_TEMPR18[0] }), .DB_DETECT( int_DB_DETECT_NG[18] ), .SB_CORRECT(int_SB_CORRECT_NG[18] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[18] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[4] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[4] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[10]  (.A(CFG3_14_Y), .B(
        CFG3_4_Y), .Y(\BLKX2[10] ));
    OR4 OR4_639 (.A(sel_R_DATA_TEMPR80[25] ), .B(sel_R_DATA_TEMPR81[25] ), 
        .C(sel_R_DATA_TEMPR82[25] ), .D(sel_R_DATA_TEMPR83[25] ), .Y(
        OR4_639_Y));
    OR4 OR4_1001 (.A(sel_R_DATA_TEMPR124[20] ), .B(sel_R_DATA_TEMPR125[20] ), 
        .C(sel_R_DATA_TEMPR126[20] ), .D(sel_R_DATA_TEMPR127[20] ), .Y(
        OR4_1001_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%15%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R15C0 (.A_DOUT({
        nc480, nc481, nc482, nc483, nc484,int_R_DATA_TEMPR15[31] , 
       int_R_DATA_TEMPR15[30] ,int_R_DATA_TEMPR15[29] , 
       int_R_DATA_TEMPR15[28] ,int_R_DATA_TEMPR15[27] , 
       int_R_DATA_TEMPR15[26] ,int_R_DATA_TEMPR15[25] , 
       int_R_DATA_TEMPR15[24] ,int_R_DATA_TEMPR15[23] , 
       int_R_DATA_TEMPR15[22] ,int_R_DATA_TEMPR15[21] , 
       int_R_DATA_TEMPR15[20] ,int_R_DATA_TEMPR15[19] , 
       int_R_DATA_TEMPR15[18] ,int_R_DATA_TEMPR15[17] }), .B_DOUT({nc485, 
        nc486, nc487,int_R_DATA_TEMPR15[16] ,int_R_DATA_TEMPR15[15] , 
       int_R_DATA_TEMPR15[14] ,int_R_DATA_TEMPR15[13] , 
       int_R_DATA_TEMPR15[12] ,int_R_DATA_TEMPR15[11] , 
       int_R_DATA_TEMPR15[10] ,int_R_DATA_TEMPR15[9] ,int_R_DATA_TEMPR15[8] , 
       int_R_DATA_TEMPR15[7] ,int_R_DATA_TEMPR15[6] ,int_R_DATA_TEMPR15[5] , 
       int_R_DATA_TEMPR15[4] ,int_R_DATA_TEMPR15[3] ,int_R_DATA_TEMPR15[2] , 
       int_R_DATA_TEMPR15[1] ,int_R_DATA_TEMPR15[0] }), .DB_DETECT( int_DB_DETECT_NG[15] ), .SB_CORRECT(int_SB_CORRECT_NG[15] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[15] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_345 (.A(sel_R_DATA_TEMPR44[31] ), .B(sel_R_DATA_TEMPR45[31] ), 
        .C(sel_R_DATA_TEMPR46[31] ), .D(sel_R_DATA_TEMPR47[31] ), .Y(
        OR4_345_Y));
    AND4 \AND4DB_DETECT[17]  (.A(sel_DB_DETECT_NG[17] ), .B(
        \BLKY2_pipe[4] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[17] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%57%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R57C0 (.A_DOUT({
        nc488, nc489, nc490, nc491, nc492,int_R_DATA_TEMPR57[31] , 
       int_R_DATA_TEMPR57[30] ,int_R_DATA_TEMPR57[29] , 
       int_R_DATA_TEMPR57[28] ,int_R_DATA_TEMPR57[27] , 
       int_R_DATA_TEMPR57[26] ,int_R_DATA_TEMPR57[25] , 
       int_R_DATA_TEMPR57[24] ,int_R_DATA_TEMPR57[23] , 
       int_R_DATA_TEMPR57[22] ,int_R_DATA_TEMPR57[21] , 
       int_R_DATA_TEMPR57[20] ,int_R_DATA_TEMPR57[19] , 
       int_R_DATA_TEMPR57[18] ,int_R_DATA_TEMPR57[17] }), .B_DOUT({nc493, 
        nc494, nc495,int_R_DATA_TEMPR57[16] ,int_R_DATA_TEMPR57[15] , 
       int_R_DATA_TEMPR57[14] ,int_R_DATA_TEMPR57[13] , 
       int_R_DATA_TEMPR57[12] ,int_R_DATA_TEMPR57[11] , 
       int_R_DATA_TEMPR57[10] ,int_R_DATA_TEMPR57[9] ,int_R_DATA_TEMPR57[8] , 
       int_R_DATA_TEMPR57[7] ,int_R_DATA_TEMPR57[6] ,int_R_DATA_TEMPR57[5] , 
       int_R_DATA_TEMPR57[4] ,int_R_DATA_TEMPR57[3] ,int_R_DATA_TEMPR57[2] , 
       int_R_DATA_TEMPR57[1] ,int_R_DATA_TEMPR57[0] }), .DB_DETECT( int_DB_DETECT_NG[57] ), .SB_CORRECT(int_SB_CORRECT_NG[57] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[57] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[14] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_236 (.A(sel_R_DATA_TEMPR8[5] ), .B(sel_R_DATA_TEMPR9[5] ), .C(sel_R_DATA_TEMPR10[5] ), .D(sel_R_DATA_TEMPR11[5] ), .Y(OR4_236_Y));
    OR4 OR4_1226 (.A(sel_R_DATA_TEMPR80[1] ), .B(sel_R_DATA_TEMPR81[1] ), .C(sel_R_DATA_TEMPR82[1] ), .D(sel_R_DATA_TEMPR83[1] ), .Y(OR4_1226_Y));
    AND4 \AND4SB_CORRECT[122]  (.A(sel_SB_CORRECT_NG[122] ), .B(
        \BLKY2_pipe[30] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[122] ));
    OR2 OR2_7 (.A(sel_R_DATA_TEMPR84[1] ), .B(sel_R_DATA_TEMPR85[1] ), .Y(
        OR2_7_Y));
    OR4 OR4_73 (.A(sel_R_DATA_TEMPR72[11] ), .B(sel_R_DATA_TEMPR73[11] ), .C(sel_R_DATA_TEMPR74[11] ), .D(sel_R_DATA_TEMPR75[11] ), .Y(OR4_73_Y));
    OR4 OR4_1042 (.A(OR4_1238_Y), .B(OR4_326_Y), .C(OR4_983_Y), .D(
        OR4_1224_Y), .Y(OR4_1042_Y));
    OR4 OR4_195 (.A(sel_R_DATA_TEMPR8[23] ), .B(sel_R_DATA_TEMPR9[23] ), .C(sel_R_DATA_TEMPR10[23] ), .D(sel_R_DATA_TEMPR11[23] ), .Y(OR4_195_Y));
    AND4 \AND4SB_CORRECT[62]  (.A(sel_SB_CORRECT_NG[62] ), .B(
        \BLKY2_pipe[15] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[62] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%66%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R66C0 (.A_DOUT({
        nc496, nc497, nc498, nc499, nc500,int_R_DATA_TEMPR66[31] , 
       int_R_DATA_TEMPR66[30] ,int_R_DATA_TEMPR66[29] , 
       int_R_DATA_TEMPR66[28] ,int_R_DATA_TEMPR66[27] , 
       int_R_DATA_TEMPR66[26] ,int_R_DATA_TEMPR66[25] , 
       int_R_DATA_TEMPR66[24] ,int_R_DATA_TEMPR66[23] , 
       int_R_DATA_TEMPR66[22] ,int_R_DATA_TEMPR66[21] , 
       int_R_DATA_TEMPR66[20] ,int_R_DATA_TEMPR66[19] , 
       int_R_DATA_TEMPR66[18] ,int_R_DATA_TEMPR66[17] }), .B_DOUT({nc501, 
        nc502, nc503,int_R_DATA_TEMPR66[16] ,int_R_DATA_TEMPR66[15] , 
       int_R_DATA_TEMPR66[14] ,int_R_DATA_TEMPR66[13] , 
       int_R_DATA_TEMPR66[12] ,int_R_DATA_TEMPR66[11] , 
       int_R_DATA_TEMPR66[10] ,int_R_DATA_TEMPR66[9] ,int_R_DATA_TEMPR66[8] , 
       int_R_DATA_TEMPR66[7] ,int_R_DATA_TEMPR66[6] ,int_R_DATA_TEMPR66[5] , 
       int_R_DATA_TEMPR66[4] ,int_R_DATA_TEMPR66[3] ,int_R_DATA_TEMPR66[2] , 
       int_R_DATA_TEMPR66[1] ,int_R_DATA_TEMPR66[0] }), .DB_DETECT( int_DB_DETECT_NG[66] ), .SB_CORRECT(int_SB_CORRECT_NG[66] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[66] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[16] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[16] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_252 (.A(OR4_629_Y), .B(OR2_32_Y), .C(sel_R_DATA_TEMPR86[10] ), 
        .D(sel_R_DATA_TEMPR87[10] ), .Y(OR4_252_Y));
    OR4 OR4_1090 (.A(OR4_409_Y), .B(OR4_777_Y), .C(OR4_225_Y), .D(
        OR4_489_Y), .Y(OR4_1090_Y));
    OR4 OR4_1328 (.A(sel_R_DATA_TEMPR44[23] ), .B(sel_R_DATA_TEMPR45[23] ), 
        .C(sel_R_DATA_TEMPR46[23] ), .D(sel_R_DATA_TEMPR47[23] ), .Y(
        OR4_1328_Y));
    OR4 OR4_289 (.A(sel_R_DATA_TEMPR24[19] ), .B(sel_R_DATA_TEMPR25[19] ), 
        .C(sel_R_DATA_TEMPR26[19] ), .D(sel_R_DATA_TEMPR27[19] ), .Y(
        OR4_289_Y));
    OR4 OR4_1003 (.A(OR4_498_Y), .B(OR4_347_Y), .C(OR4_1236_Y), .D(
        OR4_285_Y), .Y(OR4_1003_Y));
    OR4 OR4_907 (.A(sel_R_DATA_TEMPR56[29] ), .B(sel_R_DATA_TEMPR57[29] ), 
        .C(sel_R_DATA_TEMPR58[29] ), .D(sel_R_DATA_TEMPR59[29] ), .Y(
        OR4_907_Y));
    OR4 OR4_497 (.A(sel_R_DATA_TEMPR60[19] ), .B(sel_R_DATA_TEMPR61[19] ), 
        .C(sel_R_DATA_TEMPR62[19] ), .D(sel_R_DATA_TEMPR63[19] ), .Y(
        OR4_497_Y));
    OR2 OR2_32 (.A(sel_R_DATA_TEMPR84[10] ), .B(sel_R_DATA_TEMPR85[10] ), .Y(
        OR2_32_Y));
    OR4 OR4_634 (.A(sel_R_DATA_TEMPR36[3] ), .B(sel_R_DATA_TEMPR37[3] ), .C(sel_R_DATA_TEMPR38[3] ), .D(sel_R_DATA_TEMPR39[3] ), .Y(OR4_634_Y));
    OR4 OR4_1185 (.A(sel_R_DATA_TEMPR76[5] ), .B(sel_R_DATA_TEMPR77[5] ), .C(sel_R_DATA_TEMPR78[5] ), .D(sel_R_DATA_TEMPR79[5] ), .Y(OR4_1185_Y));
    OR2 OR2_1 (.A(sel_R_DATA_TEMPR84[4] ), .B(sel_R_DATA_TEMPR85[4] ), .Y(
        OR2_1_Y));
    OR4 OR4_464 (.A(sel_R_DATA_TEMPR36[11] ), .B(sel_R_DATA_TEMPR37[11] ), 
        .C(sel_R_DATA_TEMPR38[11] ), .D(sel_R_DATA_TEMPR39[11] ), .Y(
        OR4_464_Y));
    AND4 \AND4SB_CORRECT[58]  (.A(sel_SB_CORRECT_NG[58] ), .B(
        \BLKY2_pipe[14] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[58] ));
    OR4 OR4_977 (.A(OR4_280_Y), .B(OR4_353_Y), .C(OR4_796_Y), .D(
        OR4_1199_Y), .Y(OR4_977_Y));
    OR4 OR4_1081 (.A(sel_R_DATA_TEMPR80[4] ), .B(sel_R_DATA_TEMPR81[4] ), .C(sel_R_DATA_TEMPR82[4] ), .D(sel_R_DATA_TEMPR83[4] ), .Y(OR4_1081_Y));
    OR4 OR4_210 (.A(OR4_1348_Y), .B(OR4_339_Y), .C(OR4_1162_Y), .D(
        OR4_33_Y), .Y(OR4_210_Y));
    OR4 OR4_742 (.A(sel_R_DATA_TEMPR48[4] ), .B(sel_R_DATA_TEMPR49[4] ), .C(sel_R_DATA_TEMPR50[4] ), .D(sel_R_DATA_TEMPR51[4] ), .Y(OR4_742_Y));
    AND4 \AND4SB_CORRECT[100]  (.A(sel_SB_CORRECT_NG[100] ), .B(
        \BLKY2_pipe[25] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[100] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%2%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R2C0 (.A_DOUT({
        nc504, nc505, nc506, nc507, nc508,int_R_DATA_TEMPR2[31] , 
       int_R_DATA_TEMPR2[30] ,int_R_DATA_TEMPR2[29] ,int_R_DATA_TEMPR2[28] , 
       int_R_DATA_TEMPR2[27] ,int_R_DATA_TEMPR2[26] ,int_R_DATA_TEMPR2[25] , 
       int_R_DATA_TEMPR2[24] ,int_R_DATA_TEMPR2[23] ,int_R_DATA_TEMPR2[22] , 
       int_R_DATA_TEMPR2[21] ,int_R_DATA_TEMPR2[20] ,int_R_DATA_TEMPR2[19] , 
       int_R_DATA_TEMPR2[18] ,int_R_DATA_TEMPR2[17] }), .B_DOUT({nc509, 
        nc510, nc511,int_R_DATA_TEMPR2[16] ,int_R_DATA_TEMPR2[15] , 
       int_R_DATA_TEMPR2[14] ,int_R_DATA_TEMPR2[13] ,int_R_DATA_TEMPR2[12] , 
       int_R_DATA_TEMPR2[11] ,int_R_DATA_TEMPR2[10] ,int_R_DATA_TEMPR2[9] , 
       int_R_DATA_TEMPR2[8] ,int_R_DATA_TEMPR2[7] ,int_R_DATA_TEMPR2[6] , 
       int_R_DATA_TEMPR2[5] ,int_R_DATA_TEMPR2[4] ,int_R_DATA_TEMPR2[3] , 
       int_R_DATA_TEMPR2[2] ,int_R_DATA_TEMPR2[1] ,int_R_DATA_TEMPR2[0] }), 
        .DB_DETECT(int_DB_DETECT_NG[2] ), .SB_CORRECT( int_SB_CORRECT_NG[2] ), .ACCESS_BUSY(\ACCESS_BUSY[2] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[0] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_517 (.A(sel_R_DATA_TEMPR40[28] ), .B(sel_R_DATA_TEMPR41[28] ), 
        .C(sel_R_DATA_TEMPR42[28] ), .D(sel_R_DATA_TEMPR43[28] ), .Y(
        OR4_517_Y));
    OR4 OR4_350 (.A(sel_R_DATA_TEMPR92[23] ), .B(sel_R_DATA_TEMPR93[23] ), 
        .C(sel_R_DATA_TEMPR94[23] ), .D(sel_R_DATA_TEMPR95[23] ), .Y(
        OR4_350_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[1]  (.A(CFG3_8_Y), .B(CFG3_12_Y)
        , .Y(\BLKX2[1] ));
    OR4 OR4_366 (.A(sel_R_DATA_TEMPR44[7] ), .B(sel_R_DATA_TEMPR45[7] ), .C(sel_R_DATA_TEMPR46[7] ), .D(sel_R_DATA_TEMPR47[7] ), .Y(OR4_366_Y));
    OR4 OR4_295 (.A(sel_R_DATA_TEMPR112[22] ), .B(sel_R_DATA_TEMPR113[22] ), 
        .C(sel_R_DATA_TEMPR114[22] ), .D(sel_R_DATA_TEMPR115[22] ), .Y(
        OR4_295_Y));
    OR4 OR4_946 (.A(OR4_1056_Y), .B(OR4_1323_Y), .C(OR4_843_Y), .D(
        OR4_192_Y), .Y(OR4_946_Y));
    OR4 OR4_1154 (.A(sel_R_DATA_TEMPR88[20] ), .B(sel_R_DATA_TEMPR89[20] ), 
        .C(sel_R_DATA_TEMPR90[20] ), .D(sel_R_DATA_TEMPR91[20] ), .Y(
        OR4_1154_Y));
    OR4 OR4_889 (.A(sel_R_DATA_TEMPR56[9] ), .B(sel_R_DATA_TEMPR57[9] ), .C(sel_R_DATA_TEMPR58[9] ), .D(sel_R_DATA_TEMPR59[9] ), .Y(OR4_889_Y));
    AND4 \AND4SB_CORRECT[13]  (.A(sel_SB_CORRECT_NG[13] ), .B(
        \BLKY2_pipe[3] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[13] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[17]  (.A(CFG3_15_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[17] ));
    OR4 OR4_892 (.A(sel_R_DATA_TEMPR4[26] ), .B(sel_R_DATA_TEMPR5[26] ), .C(sel_R_DATA_TEMPR6[26] ), .D(sel_R_DATA_TEMPR7[26] ), .Y(OR4_892_Y));
    OR4 OR4_1029 (.A(sel_R_DATA_TEMPR96[24] ), .B(sel_R_DATA_TEMPR97[24] ), 
        .C(sel_R_DATA_TEMPR98[24] ), .D(sel_R_DATA_TEMPR99[24] ), .Y(
        OR4_1029_Y));
    OR4 OR4_645 (.A(sel_R_DATA_TEMPR116[16] ), .B(sel_R_DATA_TEMPR117[16] ), 
        .C(sel_R_DATA_TEMPR118[16] ), .D(sel_R_DATA_TEMPR119[16] ), .Y(
        OR4_645_Y));
    OR4 OR4_619 (.A(sel_R_DATA_TEMPR92[0] ), .B(sel_R_DATA_TEMPR93[0] ), .C(sel_R_DATA_TEMPR94[0] ), .D(sel_R_DATA_TEMPR95[0] ), .Y(OR4_619_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[18]  (.A(CFG3_14_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[18] ));
    OR4 OR4_1110 (.A(sel_R_DATA_TEMPR24[12] ), .B(sel_R_DATA_TEMPR25[12] ), 
        .C(sel_R_DATA_TEMPR26[12] ), .D(sel_R_DATA_TEMPR27[12] ), .Y(
        OR4_1110_Y));
    OR4 OR4_853 (.A(sel_R_DATA_TEMPR112[2] ), .B(sel_R_DATA_TEMPR113[2] ), 
        .C(sel_R_DATA_TEMPR114[2] ), .D(sel_R_DATA_TEMPR115[2] ), .Y(
        OR4_853_Y));
    AND4 \AND4DB_DETECT[35]  (.A(sel_DB_DETECT_NG[35] ), .B(
        \BLKY2_pipe[8] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[35] ));
    OR4 OR4_1083 (.A(sel_R_DATA_TEMPR116[2] ), .B(sel_R_DATA_TEMPR117[2] ), 
        .C(sel_R_DATA_TEMPR118[2] ), .D(sel_R_DATA_TEMPR119[2] ), .Y(
        OR4_1083_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[13]  (.A(CFG3_22_Y), .B(
        CFG3_4_Y), .Y(\BLKX2[13] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%34%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R34C0 (.A_DOUT({
        nc512, nc513, nc514, nc515, nc516,int_R_DATA_TEMPR34[31] , 
       int_R_DATA_TEMPR34[30] ,int_R_DATA_TEMPR34[29] , 
       int_R_DATA_TEMPR34[28] ,int_R_DATA_TEMPR34[27] , 
       int_R_DATA_TEMPR34[26] ,int_R_DATA_TEMPR34[25] , 
       int_R_DATA_TEMPR34[24] ,int_R_DATA_TEMPR34[23] , 
       int_R_DATA_TEMPR34[22] ,int_R_DATA_TEMPR34[21] , 
       int_R_DATA_TEMPR34[20] ,int_R_DATA_TEMPR34[19] , 
       int_R_DATA_TEMPR34[18] ,int_R_DATA_TEMPR34[17] }), .B_DOUT({nc517, 
        nc518, nc519,int_R_DATA_TEMPR34[16] ,int_R_DATA_TEMPR34[15] , 
       int_R_DATA_TEMPR34[14] ,int_R_DATA_TEMPR34[13] , 
       int_R_DATA_TEMPR34[12] ,int_R_DATA_TEMPR34[11] , 
       int_R_DATA_TEMPR34[10] ,int_R_DATA_TEMPR34[9] ,int_R_DATA_TEMPR34[8] , 
       int_R_DATA_TEMPR34[7] ,int_R_DATA_TEMPR34[6] ,int_R_DATA_TEMPR34[5] , 
       int_R_DATA_TEMPR34[4] ,int_R_DATA_TEMPR34[3] ,int_R_DATA_TEMPR34[2] , 
       int_R_DATA_TEMPR34[1] ,int_R_DATA_TEMPR34[0] }), .DB_DETECT( int_DB_DETECT_NG[34] ), .SB_CORRECT(int_SB_CORRECT_NG[34] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[34] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[8] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[8] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4SB_CORRECT[81]  (.A(sel_SB_CORRECT_NG[81] ), .B(
        \BLKY2_pipe[20] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[81] ));
    OR4 OR4_35 (.A(sel_R_DATA_TEMPR72[17] ), .B(sel_R_DATA_TEMPR73[17] ), .C(sel_R_DATA_TEMPR74[17] ), .D(sel_R_DATA_TEMPR75[17] ), .Y(OR4_35_Y));
    OR4 OR4_1161 (.A(\DB_DETECT[44] ), .B(\DB_DETECT[45] ), .C(
        \DB_DETECT[46] ), .D(\DB_DETECT[47] ), .Y(OR4_1161_Y));
    OR4 OR4_405 (.A(sel_R_DATA_TEMPR80[23] ), .B(sel_R_DATA_TEMPR81[23] ), 
        .C(sel_R_DATA_TEMPR82[23] ), .D(sel_R_DATA_TEMPR83[23] ), .Y(
        OR4_405_Y));
    OR4 OR4_216 (.A(OR4_1318_Y), .B(OR4_1093_Y), .C(OR4_844_Y), .D(
        OR4_948_Y), .Y(OR4_216_Y));
    AND4 \AND4DB_DETECT[48]  (.A(sel_DB_DETECT_NG[48] ), .B(
        \BLKY2_pipe[12] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[48] ));
    AND4 \AND4DB_DETECT[56]  (.A(sel_DB_DETECT_NG[56] ), .B(
        \BLKY2_pipe[14] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[56] ));
    OR4 OR4_71 (.A(OR4_1350_Y), .B(OR4_1041_Y), .C(OR4_1363_Y), .D(
        OR4_586_Y), .Y(OR4_71_Y));
    AND4 \AND4DB_DETECT[51]  (.A(sel_DB_DETECT_NG[51] ), .B(
        \BLKY2_pipe[12] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[51] ));
    OR4 OR4_1258 (.A(sel_R_DATA_TEMPR68[1] ), .B(sel_R_DATA_TEMPR69[1] ), .C(sel_R_DATA_TEMPR70[1] ), .D(sel_R_DATA_TEMPR71[1] ), .Y(OR4_1258_Y));
    OR4 OR4_475 (.A(sel_R_DATA_TEMPR124[9] ), .B(sel_R_DATA_TEMPR125[9] ), 
        .C(sel_R_DATA_TEMPR126[9] ), .D(sel_R_DATA_TEMPR127[9] ), .Y(
        OR4_475_Y));
    OR4 OR4_125 (.A(sel_R_DATA_TEMPR92[30] ), .B(sel_R_DATA_TEMPR93[30] ), 
        .C(sel_R_DATA_TEMPR94[30] ), .D(sel_R_DATA_TEMPR95[30] ), .Y(
        OR4_125_Y));
    OR4 OR4_493 (.A(sel_R_DATA_TEMPR96[9] ), .B(sel_R_DATA_TEMPR97[9] ), .C(sel_R_DATA_TEMPR98[9] ), .D(sel_R_DATA_TEMPR99[9] ), .Y(OR4_493_Y));
    OR4 OR4_1137 (.A(sel_R_DATA_TEMPR68[20] ), .B(sel_R_DATA_TEMPR69[20] ), 
        .C(sel_R_DATA_TEMPR70[20] ), .D(sel_R_DATA_TEMPR71[20] ), .Y(
        OR4_1137_Y));
    OR4 OR4_691 (.A(sel_R_DATA_TEMPR100[17] ), .B(sel_R_DATA_TEMPR101[17] ), 
        .C(sel_R_DATA_TEMPR102[17] ), .D(sel_R_DATA_TEMPR103[17] ), .Y(
        OR4_691_Y));
    OR4 OR4_614 (.A(sel_R_DATA_TEMPR24[15] ), .B(sel_R_DATA_TEMPR25[15] ), 
        .C(sel_R_DATA_TEMPR26[15] ), .D(sel_R_DATA_TEMPR27[15] ), .Y(
        OR4_614_Y));
    AND4 \AND4SB_CORRECT[14]  (.A(sel_SB_CORRECT_NG[14] ), .B(
        \BLKY2_pipe[3] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[14] ));
    OR4 OR4_427 (.A(OR4_770_Y), .B(OR4_114_Y), .C(OR4_789_Y), .D(
        OR4_1014_Y), .Y(OR4_427_Y));
    OR4 OR4_1008 (.A(OR4_371_Y), .B(OR4_914_Y), .C(OR4_1376_Y), .D(
        OR4_366_Y), .Y(OR4_1008_Y));
    OR4 OR4_787 (.A(OR4_493_Y), .B(OR4_743_Y), .C(OR4_290_Y), .D(
        OR4_999_Y), .Y(OR4_787_Y));
    OR4 OR4_298 (.A(OR4_967_Y), .B(OR4_470_Y), .C(OR4_665_Y), .D(
        OR4_1165_Y), .Y(OR4_298_Y));
    OR4 \OR4_R_DATA[27]  (.A(OR4_176_Y), .B(OR4_831_Y), .C(OR4_1203_Y), 
        .D(OR4_1327_Y), .Y(R_DATA[27]));
    OR4 OR4_784 (.A(sel_R_DATA_TEMPR64[30] ), .B(sel_R_DATA_TEMPR65[30] ), 
        .C(sel_R_DATA_TEMPR66[30] ), .D(sel_R_DATA_TEMPR67[30] ), .Y(
        OR4_784_Y));
    AND4 \AND4DB_DETECT[27]  (.A(sel_DB_DETECT_NG[27] ), .B(
        \BLKY2_pipe[6] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[27] ));
    OR4 OR4_1310 (.A(OR4_149_Y), .B(OR4_637_Y), .C(OR4_1309_Y), .D(
        OR4_137_Y), .Y(OR4_1310_Y));
    AND4 \AND4SB_CORRECT[121]  (.A(sel_SB_CORRECT_NG[121] ), .B(
        \BLKY2_pipe[30] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[121] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%40%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R40C0 (.A_DOUT({
        nc520, nc521, nc522, nc523, nc524,int_R_DATA_TEMPR40[31] , 
       int_R_DATA_TEMPR40[30] ,int_R_DATA_TEMPR40[29] , 
       int_R_DATA_TEMPR40[28] ,int_R_DATA_TEMPR40[27] , 
       int_R_DATA_TEMPR40[26] ,int_R_DATA_TEMPR40[25] , 
       int_R_DATA_TEMPR40[24] ,int_R_DATA_TEMPR40[23] , 
       int_R_DATA_TEMPR40[22] ,int_R_DATA_TEMPR40[21] , 
       int_R_DATA_TEMPR40[20] ,int_R_DATA_TEMPR40[19] , 
       int_R_DATA_TEMPR40[18] ,int_R_DATA_TEMPR40[17] }), .B_DOUT({nc525, 
        nc526, nc527,int_R_DATA_TEMPR40[16] ,int_R_DATA_TEMPR40[15] , 
       int_R_DATA_TEMPR40[14] ,int_R_DATA_TEMPR40[13] , 
       int_R_DATA_TEMPR40[12] ,int_R_DATA_TEMPR40[11] , 
       int_R_DATA_TEMPR40[10] ,int_R_DATA_TEMPR40[9] ,int_R_DATA_TEMPR40[8] , 
       int_R_DATA_TEMPR40[7] ,int_R_DATA_TEMPR40[6] ,int_R_DATA_TEMPR40[5] , 
       int_R_DATA_TEMPR40[4] ,int_R_DATA_TEMPR40[3] ,int_R_DATA_TEMPR40[2] , 
       int_R_DATA_TEMPR40[1] ,int_R_DATA_TEMPR40[0] }), .DB_DETECT( int_DB_DETECT_NG[40] ), .SB_CORRECT(int_SB_CORRECT_NG[40] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[40] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[10] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[10] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_28 (.A(sel_R_DATA_TEMPR76[11] ), .B(sel_R_DATA_TEMPR77[11] ), .C(sel_R_DATA_TEMPR78[11] ), .D(sel_R_DATA_TEMPR79[11] ), .Y(OR4_28_Y));
    OR4 OR4_1277 (.A(OR4_314_Y), .B(OR4_531_Y), .C(OR4_110_Y), .D(
        OR4_1287_Y), .Y(OR4_1277_Y));
    OR4 OR4_640 (.A(sel_R_DATA_TEMPR120[29] ), .B(sel_R_DATA_TEMPR121[29] ), 
        .C(sel_R_DATA_TEMPR122[29] ), .D(sel_R_DATA_TEMPR123[29] ), .Y(
        OR4_640_Y));
    OR4 OR4_881 (.A(OR4_681_Y), .B(OR4_1387_Y), .C(OR4_459_Y), .D(
        OR4_1328_Y), .Y(OR4_881_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%111%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R111C0 (.A_DOUT({
        nc528, nc529, nc530, nc531, nc532,int_R_DATA_TEMPR111[31] , 
       int_R_DATA_TEMPR111[30] ,int_R_DATA_TEMPR111[29] , 
       int_R_DATA_TEMPR111[28] ,int_R_DATA_TEMPR111[27] , 
       int_R_DATA_TEMPR111[26] ,int_R_DATA_TEMPR111[25] , 
       int_R_DATA_TEMPR111[24] ,int_R_DATA_TEMPR111[23] , 
       int_R_DATA_TEMPR111[22] ,int_R_DATA_TEMPR111[21] , 
       int_R_DATA_TEMPR111[20] ,int_R_DATA_TEMPR111[19] , 
       int_R_DATA_TEMPR111[18] ,int_R_DATA_TEMPR111[17] }), .B_DOUT({nc533, 
        nc534, nc535,int_R_DATA_TEMPR111[16] ,int_R_DATA_TEMPR111[15] , 
       int_R_DATA_TEMPR111[14] ,int_R_DATA_TEMPR111[13] , 
       int_R_DATA_TEMPR111[12] ,int_R_DATA_TEMPR111[11] , 
       int_R_DATA_TEMPR111[10] ,int_R_DATA_TEMPR111[9] , 
       int_R_DATA_TEMPR111[8] ,int_R_DATA_TEMPR111[7] , 
       int_R_DATA_TEMPR111[6] ,int_R_DATA_TEMPR111[5] , 
       int_R_DATA_TEMPR111[4] ,int_R_DATA_TEMPR111[3] , 
       int_R_DATA_TEMPR111[2] ,int_R_DATA_TEMPR111[1] , 
       int_R_DATA_TEMPR111[0] }), .DB_DETECT(int_DB_DETECT_NG[111] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[111] ), .ACCESS_BUSY(
        ACCESS_BUSY[111] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[27] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[27] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_164 (.A(sel_R_DATA_TEMPR80[22] ), .B(sel_R_DATA_TEMPR81[22] ), 
        .C(sel_R_DATA_TEMPR82[22] ), .D(sel_R_DATA_TEMPR83[22] ), .Y(
        OR4_164_Y));
    OR4 OR4_404 (.A(sel_R_DATA_TEMPR48[16] ), .B(sel_R_DATA_TEMPR49[16] ), 
        .C(sel_R_DATA_TEMPR50[16] ), .D(sel_R_DATA_TEMPR51[16] ), .Y(
        OR4_404_Y));
    OR4 OR4_225 (.A(sel_R_DATA_TEMPR8[0] ), .B(sel_R_DATA_TEMPR9[0] ), .C(sel_R_DATA_TEMPR10[0] ), .D(sel_R_DATA_TEMPR11[0] ), .Y(OR4_225_Y));
    OR4 OR4_555 (.A(sel_R_DATA_TEMPR64[4] ), .B(sel_R_DATA_TEMPR65[4] ), .C(sel_R_DATA_TEMPR66[4] ), .D(sel_R_DATA_TEMPR67[4] ), .Y(OR4_555_Y));
    OR4 OR4_347 (.A(sel_R_DATA_TEMPR100[30] ), .B(sel_R_DATA_TEMPR101[30] ), 
        .C(sel_R_DATA_TEMPR102[30] ), .D(sel_R_DATA_TEMPR103[30] ), .Y(
        OR4_347_Y));
    OR4 OR4_140 (.A(OR4_1143_Y), .B(OR4_993_Y), .C(OR4_1117_Y), .D(
        OR4_84_Y), .Y(OR4_140_Y));
    OR4 OR4_822 (.A(OR4_1212_Y), .B(OR4_437_Y), .C(OR4_411_Y), .D(
        OR4_1064_Y), .Y(OR4_822_Y));
    OR4 OR4_1374 (.A(sel_R_DATA_TEMPR36[30] ), .B(sel_R_DATA_TEMPR37[30] ), 
        .C(sel_R_DATA_TEMPR38[30] ), .D(sel_R_DATA_TEMPR39[30] ), .Y(
        OR4_1374_Y));
    OR4 OR4_1065 (.A(sel_R_DATA_TEMPR32[12] ), .B(sel_R_DATA_TEMPR33[12] ), 
        .C(sel_R_DATA_TEMPR34[12] ), .D(sel_R_DATA_TEMPR35[12] ), .Y(
        OR4_1065_Y));
    AND4 \AND4DB_DETECT[127]  (.A(sel_DB_DETECT_NG[127] ), .B(
        \BLKY2_pipe[31] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[127] ));
    AND4 \AND4SB_CORRECT[127]  (.A(sel_SB_CORRECT_NG[127] ), .B(
        \BLKY2_pipe[31] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[127] ));
    OR4 OR4_474 (.A(OR4_570_Y), .B(OR4_830_Y), .C(OR4_1039_Y), .D(
        OR4_870_Y), .Y(OR4_474_Y));
    OR4 OR4_1191 (.A(sel_R_DATA_TEMPR92[27] ), .B(sel_R_DATA_TEMPR93[27] ), 
        .C(sel_R_DATA_TEMPR94[27] ), .D(sel_R_DATA_TEMPR95[27] ), .Y(
        OR4_1191_Y));
    OR4 OR4_306 (.A(sel_R_DATA_TEMPR112[9] ), .B(sel_R_DATA_TEMPR113[9] ), 
        .C(sel_R_DATA_TEMPR114[9] ), .D(sel_R_DATA_TEMPR115[9] ), .Y(
        OR4_306_Y));
    OR4 OR4_1088 (.A(sel_R_DATA_TEMPR76[22] ), .B(sel_R_DATA_TEMPR77[22] ), 
        .C(sel_R_DATA_TEMPR78[22] ), .D(sel_R_DATA_TEMPR79[22] ), .Y(
        OR4_1088_Y));
    OR4 OR4_963 (.A(OR4_112_Y), .B(OR4_753_Y), .C(OR4_728_Y), .D(
        OR4_8_Y), .Y(OR4_963_Y));
    AND4 \AND4SB_CORRECT[35]  (.A(sel_SB_CORRECT_NG[35] ), .B(
        \BLKY2_pipe[8] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[35] ));
    AND4 \AND4SB_CORRECT[36]  (.A(sel_SB_CORRECT_NG[36] ), .B(
        \BLKY2_pipe[9] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[36] ));
    OR4 OR4_748 (.A(sel_R_DATA_TEMPR16[19] ), .B(sel_R_DATA_TEMPR17[19] ), 
        .C(sel_R_DATA_TEMPR18[19] ), .D(sel_R_DATA_TEMPR19[19] ), .Y(
        OR4_748_Y));
    OR4 OR4_653 (.A(OR4_70_Y), .B(OR4_1028_Y), .C(OR4_1068_Y), .D(
        OR4_203_Y), .Y(OR4_653_Y));
    OR4 OR4_1155 (.A(sel_R_DATA_TEMPR108[3] ), .B(sel_R_DATA_TEMPR109[3] ), 
        .C(sel_R_DATA_TEMPR110[3] ), .D(sel_R_DATA_TEMPR111[3] ), .Y(
        OR4_1155_Y));
    OR4 OR4_376 (.A(OR4_1257_Y), .B(OR4_991_Y), .C(OR4_965_Y), .D(
        OR4_262_Y), .Y(OR4_376_Y));
    OR4 OR4_866 (.A(OR4_523_Y), .B(OR4_774_Y), .C(OR4_318_Y), .D(
        OR4_1038_Y), .Y(OR4_866_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[18]  (.A(CFG3_0_Y), .B(CFG3_9_Y)
        , .Y(\BLKY2[18] ));
    OR4 OR4_1051 (.A(sel_R_DATA_TEMPR104[19] ), .B(sel_R_DATA_TEMPR105[19] ), 
        .C(sel_R_DATA_TEMPR106[19] ), .D(sel_R_DATA_TEMPR107[19] ), .Y(
        OR4_1051_Y));
    OR4 OR4_761 (.A(sel_R_DATA_TEMPR68[12] ), .B(sel_R_DATA_TEMPR69[12] ), 
        .C(sel_R_DATA_TEMPR70[12] ), .D(sel_R_DATA_TEMPR71[12] ), .Y(
        OR4_761_Y));
    OR4 OR4_1127 (.A(sel_R_DATA_TEMPR60[29] ), .B(sel_R_DATA_TEMPR61[29] ), 
        .C(sel_R_DATA_TEMPR62[29] ), .D(sel_R_DATA_TEMPR63[29] ), .Y(
        OR4_1127_Y));
    OR4 OR4_1215 (.A(sel_R_DATA_TEMPR36[26] ), .B(sel_R_DATA_TEMPR37[26] ), 
        .C(sel_R_DATA_TEMPR38[26] ), .D(sel_R_DATA_TEMPR39[26] ), .Y(
        OR4_1215_Y));
    AND4 \AND4SB_CORRECT[99]  (.A(sel_SB_CORRECT_NG[99] ), .B(
        \BLKY2_pipe[24] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[99] ));
    OR4 OR4_423 (.A(sel_R_DATA_TEMPR104[6] ), .B(sel_R_DATA_TEMPR105[6] ), 
        .C(sel_R_DATA_TEMPR106[6] ), .D(sel_R_DATA_TEMPR107[6] ), .Y(
        OR4_423_Y));
    OR4 OR4_621 (.A(OR4_422_Y), .B(OR4_788_Y), .C(OR4_236_Y), .D(
        OR4_500_Y), .Y(OR4_621_Y));
    OR4 OR4_84 (.A(sel_R_DATA_TEMPR124[12] ), .B(sel_R_DATA_TEMPR125[12] ), 
        .C(sel_R_DATA_TEMPR126[12] ), .D(sel_R_DATA_TEMPR127[12] ), .Y(
        OR4_84_Y));
    OR4 OR4_1230 (.A(sel_R_DATA_TEMPR48[1] ), .B(sel_R_DATA_TEMPR49[1] ), .C(sel_R_DATA_TEMPR50[1] ), .D(sel_R_DATA_TEMPR51[1] ), .Y(OR4_1230_Y));
    OR4 OR4_847 (.A(OR4_1176_Y), .B(OR4_327_Y), .C(OR4_771_Y), .D(
        OR4_278_Y), .Y(OR4_847_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[13]  (.A(CFG3_11_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[13] ));
    OR4 OR4_148 (.A(sel_R_DATA_TEMPR20[3] ), .B(sel_R_DATA_TEMPR21[3] ), .C(sel_R_DATA_TEMPR22[3] ), .D(sel_R_DATA_TEMPR23[3] ), .Y(OR4_148_Y));
    OR4 OR4_944 (.A(sel_R_DATA_TEMPR60[18] ), .B(sel_R_DATA_TEMPR61[18] ), 
        .C(sel_R_DATA_TEMPR62[18] ), .D(sel_R_DATA_TEMPR63[18] ), .Y(
        OR4_944_Y));
    OR4 OR4_228 (.A(OR4_625_Y), .B(OR4_412_Y), .C(OR4_167_Y), .D(
        OR4_481_Y), .Y(OR4_228_Y));
    OR4 OR4_838 (.A(sel_R_DATA_TEMPR44[21] ), .B(sel_R_DATA_TEMPR45[21] ), 
        .C(sel_R_DATA_TEMPR46[21] ), .D(sel_R_DATA_TEMPR47[21] ), .Y(
        OR4_838_Y));
    OR4 OR4_1379 (.A(sel_R_DATA_TEMPR4[25] ), .B(sel_R_DATA_TEMPR5[25] ), .C(sel_R_DATA_TEMPR6[25] ), .D(sel_R_DATA_TEMPR7[25] ), .Y(OR4_1379_Y));
    OR4 OR4_987 (.A(sel_R_DATA_TEMPR76[27] ), .B(sel_R_DATA_TEMPR77[27] ), 
        .C(sel_R_DATA_TEMPR78[27] ), .D(sel_R_DATA_TEMPR79[27] ), .Y(
        OR4_987_Y));
    OR4 OR4_959 (.A(sel_R_DATA_TEMPR24[8] ), .B(sel_R_DATA_TEMPR25[8] ), .C(sel_R_DATA_TEMPR26[8] ), .D(sel_R_DATA_TEMPR27[8] ), .Y(OR4_959_Y));
    OR4 OR4_950 (.A(sel_R_DATA_TEMPR0[13] ), .B(sel_R_DATA_TEMPR1[13] ), .C(sel_R_DATA_TEMPR2[13] ), .D(sel_R_DATA_TEMPR3[13] ), .Y(OR4_950_Y));
    OR4 OR4_566 (.A(sel_R_DATA_TEMPR56[11] ), .B(sel_R_DATA_TEMPR57[11] ), 
        .C(sel_R_DATA_TEMPR58[11] ), .D(sel_R_DATA_TEMPR59[11] ), .Y(
        OR4_566_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[3]  (.D(\BLKY2[3] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[3] ));
    OR4 OR4_591 (.A(OR4_1179_Y), .B(OR4_3_Y), .C(OR4_166_Y), .D(
        OR4_307_Y), .Y(OR4_591_Y));
    OR4 OR4_1053 (.A(sel_R_DATA_TEMPR100[16] ), .B(sel_R_DATA_TEMPR101[16] ), 
        .C(sel_R_DATA_TEMPR102[16] ), .D(sel_R_DATA_TEMPR103[16] ), .Y(
        OR4_1053_Y));
    CFG3 #( .INIT(8'h20) )  CFG3_4 (.A(W_EN), .B(W_ADDR[15]), .C(
        W_ADDR[14]), .Y(CFG3_4_Y));
    OR4 OR4_1070 (.A(\SB_CORRECT[92] ), .B(\SB_CORRECT[93] ), .C(
        \SB_CORRECT[94] ), .D(\SB_CORRECT[95] ), .Y(OR4_1070_Y));
    AND4 \AND4DB_DETECT[86]  (.A(sel_DB_DETECT_NG[86] ), .B(
        \BLKY2_pipe[21] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[86] ));
    AND4 \AND4SB_CORRECT[77]  (.A(sel_SB_CORRECT_NG[77] ), .B(
        \BLKY2_pipe[19] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[77] ));
    OR4 OR4_1007 (.A(sel_R_DATA_TEMPR60[27] ), .B(sel_R_DATA_TEMPR61[27] ), 
        .C(sel_R_DATA_TEMPR62[27] ), .D(sel_R_DATA_TEMPR63[27] ), .Y(
        OR4_1007_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[9]  (.A(CFG3_8_Y), .B(CFG3_4_Y), 
        .Y(\BLKX2[9] ));
    OR4 OR4_1332 (.A(OR4_360_Y), .B(OR4_741_Y), .C(OR4_178_Y), .D(
        OR4_451_Y), .Y(OR4_1332_Y));
    AND4 \AND4DB_DETECT[49]  (.A(sel_DB_DETECT_NG[49] ), .B(
        \BLKY2_pipe[12] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[49] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%56%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R56C0 (.A_DOUT({
        nc536, nc537, nc538, nc539, nc540,int_R_DATA_TEMPR56[31] , 
       int_R_DATA_TEMPR56[30] ,int_R_DATA_TEMPR56[29] , 
       int_R_DATA_TEMPR56[28] ,int_R_DATA_TEMPR56[27] , 
       int_R_DATA_TEMPR56[26] ,int_R_DATA_TEMPR56[25] , 
       int_R_DATA_TEMPR56[24] ,int_R_DATA_TEMPR56[23] , 
       int_R_DATA_TEMPR56[22] ,int_R_DATA_TEMPR56[21] , 
       int_R_DATA_TEMPR56[20] ,int_R_DATA_TEMPR56[19] , 
       int_R_DATA_TEMPR56[18] ,int_R_DATA_TEMPR56[17] }), .B_DOUT({nc541, 
        nc542, nc543,int_R_DATA_TEMPR56[16] ,int_R_DATA_TEMPR56[15] , 
       int_R_DATA_TEMPR56[14] ,int_R_DATA_TEMPR56[13] , 
       int_R_DATA_TEMPR56[12] ,int_R_DATA_TEMPR56[11] , 
       int_R_DATA_TEMPR56[10] ,int_R_DATA_TEMPR56[9] ,int_R_DATA_TEMPR56[8] , 
       int_R_DATA_TEMPR56[7] ,int_R_DATA_TEMPR56[6] ,int_R_DATA_TEMPR56[5] , 
       int_R_DATA_TEMPR56[4] ,int_R_DATA_TEMPR56[3] ,int_R_DATA_TEMPR56[2] , 
       int_R_DATA_TEMPR56[1] ,int_R_DATA_TEMPR56[0] }), .DB_DETECT( int_DB_DETECT_NG[56] ), .SB_CORRECT(int_SB_CORRECT_NG[56] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[56] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[14] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[14] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4DB_DETECT[81]  (.A(sel_DB_DETECT_NG[81] ), .B(
        \BLKY2_pipe[20] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[81] ));
    OR4 OR4_153 (.A(sel_R_DATA_TEMPR8[16] ), .B(sel_R_DATA_TEMPR9[16] ), .C(sel_R_DATA_TEMPR10[16] ), .D(sel_R_DATA_TEMPR11[16] ), .Y(OR4_153_Y));
    OR4 OR4_1232 (.A(sel_R_DATA_TEMPR104[1] ), .B(sel_R_DATA_TEMPR105[1] ), 
        .C(sel_R_DATA_TEMPR106[1] ), .D(sel_R_DATA_TEMPR107[1] ), .Y(
        OR4_1232_Y));
    OR4 OR4_1095 (.A(sel_R_DATA_TEMPR16[15] ), .B(sel_R_DATA_TEMPR17[15] ), 
        .C(sel_R_DATA_TEMPR18[15] ), .D(sel_R_DATA_TEMPR19[15] ), .Y(
        OR4_1095_Y));
    OR4 OR4_9 (.A(OR4_335_Y), .B(OR4_1148_Y), .C(OR4_1123_Y), .D(
        OR4_399_Y), .Y(OR4_9_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[23]  (.D(\BLKY2[23] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[23] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%30%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R30C0 (.A_DOUT({
        nc544, nc545, nc546, nc547, nc548,int_R_DATA_TEMPR30[31] , 
       int_R_DATA_TEMPR30[30] ,int_R_DATA_TEMPR30[29] , 
       int_R_DATA_TEMPR30[28] ,int_R_DATA_TEMPR30[27] , 
       int_R_DATA_TEMPR30[26] ,int_R_DATA_TEMPR30[25] , 
       int_R_DATA_TEMPR30[24] ,int_R_DATA_TEMPR30[23] , 
       int_R_DATA_TEMPR30[22] ,int_R_DATA_TEMPR30[21] , 
       int_R_DATA_TEMPR30[20] ,int_R_DATA_TEMPR30[19] , 
       int_R_DATA_TEMPR30[18] ,int_R_DATA_TEMPR30[17] }), .B_DOUT({nc549, 
        nc550, nc551,int_R_DATA_TEMPR30[16] ,int_R_DATA_TEMPR30[15] , 
       int_R_DATA_TEMPR30[14] ,int_R_DATA_TEMPR30[13] , 
       int_R_DATA_TEMPR30[12] ,int_R_DATA_TEMPR30[11] , 
       int_R_DATA_TEMPR30[10] ,int_R_DATA_TEMPR30[9] ,int_R_DATA_TEMPR30[8] , 
       int_R_DATA_TEMPR30[7] ,int_R_DATA_TEMPR30[6] ,int_R_DATA_TEMPR30[5] , 
       int_R_DATA_TEMPR30[4] ,int_R_DATA_TEMPR30[3] ,int_R_DATA_TEMPR30[2] , 
       int_R_DATA_TEMPR30[1] ,int_R_DATA_TEMPR30[0] }), .DB_DETECT( int_DB_DETECT_NG[30] ), .SB_CORRECT(int_SB_CORRECT_NG[30] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[30] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[7] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_231 (.A(sel_R_DATA_TEMPR80[0] ), .B(sel_R_DATA_TEMPR81[0] ), .C(sel_R_DATA_TEMPR82[0] ), .D(sel_R_DATA_TEMPR83[0] ), .Y(OR4_231_Y));
    OR4 OR4_104 (.A(sel_R_DATA_TEMPR40[15] ), .B(sel_R_DATA_TEMPR41[15] ), 
        .C(sel_R_DATA_TEMPR42[15] ), .D(sel_R_DATA_TEMPR43[15] ), .Y(
        OR4_104_Y));
    OR4 OR4_292 (.A(sel_R_DATA_TEMPR8[19] ), .B(sel_R_DATA_TEMPR9[19] ), .C(sel_R_DATA_TEMPR10[19] ), .D(sel_R_DATA_TEMPR11[19] ), .Y(OR4_292_Y));
    OR4 OR4_DB_DETECT (.A(OR4_1392_Y), .B(OR4_109_Y), .C(OR4_592_Y), 
        .D(OR4_1249_Y), .Y(DB_DETECT));
    CFG3 #( .INIT(8'h40) )  CFG3_5 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_5_Y));
    OR4 OR4_1160 (.A(sel_R_DATA_TEMPR104[4] ), .B(sel_R_DATA_TEMPR105[4] ), 
        .C(sel_R_DATA_TEMPR106[4] ), .D(sel_R_DATA_TEMPR107[4] ), .Y(
        OR4_1160_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%74%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R74C0 (.A_DOUT({
        nc552, nc553, nc554, nc555, nc556,int_R_DATA_TEMPR74[31] , 
       int_R_DATA_TEMPR74[30] ,int_R_DATA_TEMPR74[29] , 
       int_R_DATA_TEMPR74[28] ,int_R_DATA_TEMPR74[27] , 
       int_R_DATA_TEMPR74[26] ,int_R_DATA_TEMPR74[25] , 
       int_R_DATA_TEMPR74[24] ,int_R_DATA_TEMPR74[23] , 
       int_R_DATA_TEMPR74[22] ,int_R_DATA_TEMPR74[21] , 
       int_R_DATA_TEMPR74[20] ,int_R_DATA_TEMPR74[19] , 
       int_R_DATA_TEMPR74[18] ,int_R_DATA_TEMPR74[17] }), .B_DOUT({nc557, 
        nc558, nc559,int_R_DATA_TEMPR74[16] ,int_R_DATA_TEMPR74[15] , 
       int_R_DATA_TEMPR74[14] ,int_R_DATA_TEMPR74[13] , 
       int_R_DATA_TEMPR74[12] ,int_R_DATA_TEMPR74[11] , 
       int_R_DATA_TEMPR74[10] ,int_R_DATA_TEMPR74[9] ,int_R_DATA_TEMPR74[8] , 
       int_R_DATA_TEMPR74[7] ,int_R_DATA_TEMPR74[6] ,int_R_DATA_TEMPR74[5] , 
       int_R_DATA_TEMPR74[4] ,int_R_DATA_TEMPR74[3] ,int_R_DATA_TEMPR74[2] , 
       int_R_DATA_TEMPR74[1] ,int_R_DATA_TEMPR74[0] }), .DB_DETECT( int_DB_DETECT_NG[74] ), .SB_CORRECT(int_SB_CORRECT_NG[74] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[74] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[18] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[18] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1234 (.A(sel_R_DATA_TEMPR60[30] ), .B(sel_R_DATA_TEMPR61[30] ), 
        .C(sel_R_DATA_TEMPR62[30] ), .D(sel_R_DATA_TEMPR63[30] ), .Y(
        OR4_1234_Y));
    OR4 OR4_174 (.A(\SB_CORRECT[32] ), .B(\SB_CORRECT[33] ), .C(
        \SB_CORRECT[34] ), .D(\SB_CORRECT[35] ), .Y(OR4_174_Y));
    OR4 OR4_485 (.A(OR4_1331_Y), .B(OR4_319_Y), .C(OR4_304_Y), .D(
        OR4_952_Y), .Y(OR4_485_Y));
    OR4 OR4_1337 (.A(sel_R_DATA_TEMPR76[23] ), .B(sel_R_DATA_TEMPR77[23] ), 
        .C(sel_R_DATA_TEMPR78[23] ), .D(sel_R_DATA_TEMPR79[23] ), .Y(
        OR4_1337_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[29]  (.A(CFG3_22_Y), .B(
        CFG3_7_Y), .Y(\BLKX2[29] ));
    OR4 OR4_1087 (.A(sel_R_DATA_TEMPR92[5] ), .B(sel_R_DATA_TEMPR93[5] ), .C(sel_R_DATA_TEMPR94[5] ), .D(sel_R_DATA_TEMPR95[5] ), .Y(OR4_1087_Y));
    OR4 OR4_903 (.A(sel_R_DATA_TEMPR52[18] ), .B(sel_R_DATA_TEMPR53[18] ), 
        .C(sel_R_DATA_TEMPR54[18] ), .D(sel_R_DATA_TEMPR55[18] ), .Y(
        OR4_903_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%127%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R127C0 (.A_DOUT({
        nc560, nc561, nc562, nc563, nc564,int_R_DATA_TEMPR127[31] , 
       int_R_DATA_TEMPR127[30] ,int_R_DATA_TEMPR127[29] , 
       int_R_DATA_TEMPR127[28] ,int_R_DATA_TEMPR127[27] , 
       int_R_DATA_TEMPR127[26] ,int_R_DATA_TEMPR127[25] , 
       int_R_DATA_TEMPR127[24] ,int_R_DATA_TEMPR127[23] , 
       int_R_DATA_TEMPR127[22] ,int_R_DATA_TEMPR127[21] , 
       int_R_DATA_TEMPR127[20] ,int_R_DATA_TEMPR127[19] , 
       int_R_DATA_TEMPR127[18] ,int_R_DATA_TEMPR127[17] }), .B_DOUT({nc565, 
        nc566, nc567,int_R_DATA_TEMPR127[16] ,int_R_DATA_TEMPR127[15] , 
       int_R_DATA_TEMPR127[14] ,int_R_DATA_TEMPR127[13] , 
       int_R_DATA_TEMPR127[12] ,int_R_DATA_TEMPR127[11] , 
       int_R_DATA_TEMPR127[10] ,int_R_DATA_TEMPR127[9] , 
       int_R_DATA_TEMPR127[8] ,int_R_DATA_TEMPR127[7] , 
       int_R_DATA_TEMPR127[6] ,int_R_DATA_TEMPR127[5] , 
       int_R_DATA_TEMPR127[4] ,int_R_DATA_TEMPR127[3] , 
       int_R_DATA_TEMPR127[2] ,int_R_DATA_TEMPR127[1] , 
       int_R_DATA_TEMPR127[0] }), .DB_DETECT(int_DB_DETECT_NG[127] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[127] ), .ACCESS_BUSY(
        ACCESS_BUSY[127] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[31] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[31] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4SB_CORRECT[21]  (.A(sel_SB_CORRECT_NG[21] ), .B(
        \BLKY2_pipe[5] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[21] ));
    OR4 OR4_568 (.A(sel_R_DATA_TEMPR60[14] ), .B(sel_R_DATA_TEMPR61[14] ), 
        .C(sel_R_DATA_TEMPR62[14] ), .D(sel_R_DATA_TEMPR63[14] ), .Y(
        OR4_568_Y));
    OR4 OR4_1220 (.A(sel_R_DATA_TEMPR80[29] ), .B(sel_R_DATA_TEMPR81[29] ), 
        .C(sel_R_DATA_TEMPR82[29] ), .D(sel_R_DATA_TEMPR83[29] ), .Y(
        OR4_1220_Y));
    OR4 OR4_532 (.A(sel_R_DATA_TEMPR16[9] ), .B(sel_R_DATA_TEMPR17[9] ), .C(sel_R_DATA_TEMPR18[9] ), .D(sel_R_DATA_TEMPR19[9] ), .Y(OR4_532_Y));
    OR4 OR4_56 (.A(sel_R_DATA_TEMPR64[22] ), .B(sel_R_DATA_TEMPR65[22] ), .C(sel_R_DATA_TEMPR66[22] ), .D(sel_R_DATA_TEMPR67[22] ), .Y(OR4_56_Y));
    AND4 \AND4SB_CORRECT[116]  (.A(sel_SB_CORRECT_NG[116] ), .B(
        \BLKY2_pipe[29] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[116] ));
    OR4 OR4_390 (.A(sel_R_DATA_TEMPR92[31] ), .B(sel_R_DATA_TEMPR93[31] ), 
        .C(sel_R_DATA_TEMPR94[31] ), .D(sel_R_DATA_TEMPR95[31] ), .Y(
        OR4_390_Y));
    OR4 OR4_818 (.A(sel_R_DATA_TEMPR56[21] ), .B(sel_R_DATA_TEMPR57[21] ), 
        .C(sel_R_DATA_TEMPR58[21] ), .D(sel_R_DATA_TEMPR59[21] ), .Y(
        OR4_818_Y));
    OR4 OR4_973 (.A(sel_R_DATA_TEMPR124[15] ), .B(sel_R_DATA_TEMPR125[15] ), 
        .C(sel_R_DATA_TEMPR126[15] ), .D(sel_R_DATA_TEMPR127[15] ), .Y(
        OR4_973_Y));
    OR4 OR4_806 (.A(OR4_1054_Y), .B(OR4_161_Y), .C(OR4_818_Y), .D(
        OR4_1043_Y), .Y(OR4_806_Y));
    OR4 OR4_701 (.A(sel_R_DATA_TEMPR40[20] ), .B(sel_R_DATA_TEMPR41[20] ), 
        .C(sel_R_DATA_TEMPR42[20] ), .D(sel_R_DATA_TEMPR43[20] ), .Y(
        OR4_701_Y));
    AND4 \AND4SB_CORRECT[113]  (.A(sel_SB_CORRECT_NG[113] ), .B(
        \BLKY2_pipe[28] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[113] ));
    AND4 \AND4SB_CORRECT[124]  (.A(sel_SB_CORRECT_NG[124] ), .B(
        \BLKY2_pipe[31] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[124] ));
    OR4 \OR4_R_DATA[2]  (.A(OR4_752_Y), .B(OR4_679_Y), .C(OR4_946_Y), 
        .D(OR4_1046_Y), .Y(R_DATA[2]));
    OR4 OR4_850 (.A(sel_R_DATA_TEMPR120[30] ), .B(sel_R_DATA_TEMPR121[30] ), 
        .C(sel_R_DATA_TEMPR122[30] ), .D(sel_R_DATA_TEMPR123[30] ), .Y(
        OR4_850_Y));
    AND4 \AND4SB_CORRECT[57]  (.A(sel_SB_CORRECT_NG[57] ), .B(
        \BLKY2_pipe[14] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[57] ));
    OR4 OR4_521 (.A(sel_R_DATA_TEMPR124[22] ), .B(sel_R_DATA_TEMPR125[22] ), 
        .C(sel_R_DATA_TEMPR126[22] ), .D(sel_R_DATA_TEMPR127[22] ), .Y(
        OR4_521_Y));
    OR4 OR4_1322 (.A(sel_R_DATA_TEMPR28[6] ), .B(sel_R_DATA_TEMPR29[6] ), .C(sel_R_DATA_TEMPR30[6] ), .D(sel_R_DATA_TEMPR31[6] ), .Y(OR4_1322_Y));
    OR4 OR4_876 (.A(sel_R_DATA_TEMPR92[10] ), .B(sel_R_DATA_TEMPR93[10] ), 
        .C(sel_R_DATA_TEMPR94[10] ), .D(sel_R_DATA_TEMPR95[10] ), .Y(
        OR4_876_Y));
    OR4 OR4_1058 (.A(\SB_CORRECT[52] ), .B(\SB_CORRECT[53] ), .C(
        \SB_CORRECT[54] ), .D(\SB_CORRECT[55] ), .Y(OR4_1058_Y));
    OR4 OR4_771 (.A(sel_R_DATA_TEMPR40[22] ), .B(sel_R_DATA_TEMPR41[22] ), 
        .C(sel_R_DATA_TEMPR42[22] ), .D(sel_R_DATA_TEMPR43[22] ), .Y(
        OR4_771_Y));
    OR4 OR4_152 (.A(sel_R_DATA_TEMPR0[29] ), .B(sel_R_DATA_TEMPR1[29] ), .C(sel_R_DATA_TEMPR2[29] ), .D(sel_R_DATA_TEMPR3[29] ), .Y(OR4_152_Y));
    OR4 OR4_893 (.A(OR4_622_Y), .B(OR4_468_Y), .C(OR4_151_Y), .D(
        OR4_11_Y), .Y(OR4_893_Y));
    OR4 OR4_1222 (.A(sel_R_DATA_TEMPR120[22] ), .B(sel_R_DATA_TEMPR121[22] ), 
        .C(sel_R_DATA_TEMPR122[22] ), .D(sel_R_DATA_TEMPR123[22] ), .Y(
        OR4_1222_Y));
    OR4 OR4_1360 (.A(sel_R_DATA_TEMPR124[5] ), .B(sel_R_DATA_TEMPR125[5] ), 
        .C(sel_R_DATA_TEMPR126[5] ), .D(sel_R_DATA_TEMPR127[5] ), .Y(
        OR4_1360_Y));
    OR4 OR4_466 (.A(sel_R_DATA_TEMPR28[26] ), .B(sel_R_DATA_TEMPR29[26] ), 
        .C(sel_R_DATA_TEMPR30[26] ), .D(sel_R_DATA_TEMPR31[26] ), .Y(
        OR4_466_Y));
    OR4 OR4_955 (.A(sel_R_DATA_TEMPR112[27] ), .B(sel_R_DATA_TEMPR113[27] ), 
        .C(sel_R_DATA_TEMPR114[27] ), .D(sel_R_DATA_TEMPR115[27] ), .Y(
        OR4_955_Y));
    OR4 OR4_39 (.A(sel_R_DATA_TEMPR124[25] ), .B(sel_R_DATA_TEMPR125[25] ), 
        .C(sel_R_DATA_TEMPR126[25] ), .D(sel_R_DATA_TEMPR127[25] ), .Y(
        OR4_39_Y));
    OR4 OR4_534 (.A(\DB_DETECT[100] ), .B(\DB_DETECT[101] ), .C(
        \DB_DETECT[102] ), .D(\DB_DETECT[103] ), .Y(OR4_534_Y));
    OR4 OR4_506 (.A(sel_R_DATA_TEMPR68[18] ), .B(sel_R_DATA_TEMPR69[18] ), 
        .C(sel_R_DATA_TEMPR70[18] ), .D(sel_R_DATA_TEMPR71[18] ), .Y(
        OR4_506_Y));
    OR4 OR4_211 (.A(sel_R_DATA_TEMPR100[21] ), .B(sel_R_DATA_TEMPR101[21] ), 
        .C(sel_R_DATA_TEMPR102[21] ), .D(sel_R_DATA_TEMPR103[21] ), .Y(
        OR4_211_Y));
    OR4 OR4_932 (.A(sel_R_DATA_TEMPR16[20] ), .B(sel_R_DATA_TEMPR17[20] ), 
        .C(sel_R_DATA_TEMPR18[20] ), .D(sel_R_DATA_TEMPR19[20] ), .Y(
        OR4_932_Y));
    OR4 OR4_484 (.A(sel_R_DATA_TEMPR88[11] ), .B(sel_R_DATA_TEMPR89[11] ), 
        .C(sel_R_DATA_TEMPR90[11] ), .D(sel_R_DATA_TEMPR91[11] ), .Y(
        OR4_484_Y));
    OR2 OR2_9 (.A(sel_R_DATA_TEMPR84[15] ), .B(sel_R_DATA_TEMPR85[15] ), .Y(
        OR2_9_Y));
    OR4 OR4_1014 (.A(sel_R_DATA_TEMPR28[2] ), .B(sel_R_DATA_TEMPR29[2] ), .C(sel_R_DATA_TEMPR30[2] ), .D(sel_R_DATA_TEMPR31[2] ), .Y(OR4_1014_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[22]  (.D(\BLKY2[22] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[22] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%29%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R29C0 (.A_DOUT({
        nc568, nc569, nc570, nc571, nc572,int_R_DATA_TEMPR29[31] , 
       int_R_DATA_TEMPR29[30] ,int_R_DATA_TEMPR29[29] , 
       int_R_DATA_TEMPR29[28] ,int_R_DATA_TEMPR29[27] , 
       int_R_DATA_TEMPR29[26] ,int_R_DATA_TEMPR29[25] , 
       int_R_DATA_TEMPR29[24] ,int_R_DATA_TEMPR29[23] , 
       int_R_DATA_TEMPR29[22] ,int_R_DATA_TEMPR29[21] , 
       int_R_DATA_TEMPR29[20] ,int_R_DATA_TEMPR29[19] , 
       int_R_DATA_TEMPR29[18] ,int_R_DATA_TEMPR29[17] }), .B_DOUT({nc573, 
        nc574, nc575,int_R_DATA_TEMPR29[16] ,int_R_DATA_TEMPR29[15] , 
       int_R_DATA_TEMPR29[14] ,int_R_DATA_TEMPR29[13] , 
       int_R_DATA_TEMPR29[12] ,int_R_DATA_TEMPR29[11] , 
       int_R_DATA_TEMPR29[10] ,int_R_DATA_TEMPR29[9] ,int_R_DATA_TEMPR29[8] , 
       int_R_DATA_TEMPR29[7] ,int_R_DATA_TEMPR29[6] ,int_R_DATA_TEMPR29[5] , 
       int_R_DATA_TEMPR29[4] ,int_R_DATA_TEMPR29[3] ,int_R_DATA_TEMPR29[2] , 
       int_R_DATA_TEMPR29[1] ,int_R_DATA_TEMPR29[0] }), .DB_DETECT( int_DB_DETECT_NG[29] ), .SB_CORRECT(int_SB_CORRECT_NG[29] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[29] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1190 (.A(sel_R_DATA_TEMPR44[19] ), .B(sel_R_DATA_TEMPR45[19] ), 
        .C(sel_R_DATA_TEMPR46[19] ), .D(sel_R_DATA_TEMPR47[19] ), .Y(
        OR4_1190_Y));
    OR4 OR4_576 (.A(sel_R_DATA_TEMPR28[29] ), .B(sel_R_DATA_TEMPR29[29] ), 
        .C(sel_R_DATA_TEMPR30[29] ), .D(sel_R_DATA_TEMPR31[29] ), .Y(
        OR4_576_Y));
    OR4 OR4_1224 (.A(sel_R_DATA_TEMPR60[24] ), .B(sel_R_DATA_TEMPR61[24] ), 
        .C(sel_R_DATA_TEMPR62[24] ), .D(sel_R_DATA_TEMPR63[24] ), .Y(
        OR4_1224_Y));
    AND4 \AND4SB_CORRECT[61]  (.A(sel_SB_CORRECT_NG[61] ), .B(
        \BLKY2_pipe[15] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[61] ));
    OR4 OR4_145 (.A(OR4_939_Y), .B(OR4_615_Y), .C(OR4_588_Y), .D(
        OR4_1271_Y), .Y(OR4_145_Y));
    OR4 OR4_362 (.A(sel_R_DATA_TEMPR16[4] ), .B(sel_R_DATA_TEMPR17[4] ), .C(sel_R_DATA_TEMPR18[4] ), .D(sel_R_DATA_TEMPR19[4] ), .Y(OR4_362_Y));
    OR4 OR4_222 (.A(sel_R_DATA_TEMPR88[1] ), .B(sel_R_DATA_TEMPR89[1] ), .C(sel_R_DATA_TEMPR90[1] ), .D(sel_R_DATA_TEMPR91[1] ), .Y(OR4_222_Y));
    OR4 OR4_1313 (.A(sel_R_DATA_TEMPR68[17] ), .B(sel_R_DATA_TEMPR69[17] ), 
        .C(sel_R_DATA_TEMPR70[17] ), .D(sel_R_DATA_TEMPR71[17] ), .Y(
        OR4_1313_Y));
    OR4 OR4_1143 (.A(sel_R_DATA_TEMPR112[12] ), .B(sel_R_DATA_TEMPR113[12] ), 
        .C(sel_R_DATA_TEMPR114[12] ), .D(sel_R_DATA_TEMPR115[12] ), .Y(
        OR4_1143_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%68%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R68C0 (.A_DOUT({
        nc576, nc577, nc578, nc579, nc580,int_R_DATA_TEMPR68[31] , 
       int_R_DATA_TEMPR68[30] ,int_R_DATA_TEMPR68[29] , 
       int_R_DATA_TEMPR68[28] ,int_R_DATA_TEMPR68[27] , 
       int_R_DATA_TEMPR68[26] ,int_R_DATA_TEMPR68[25] , 
       int_R_DATA_TEMPR68[24] ,int_R_DATA_TEMPR68[23] , 
       int_R_DATA_TEMPR68[22] ,int_R_DATA_TEMPR68[21] , 
       int_R_DATA_TEMPR68[20] ,int_R_DATA_TEMPR68[19] , 
       int_R_DATA_TEMPR68[18] ,int_R_DATA_TEMPR68[17] }), .B_DOUT({nc581, 
        nc582, nc583,int_R_DATA_TEMPR68[16] ,int_R_DATA_TEMPR68[15] , 
       int_R_DATA_TEMPR68[14] ,int_R_DATA_TEMPR68[13] , 
       int_R_DATA_TEMPR68[12] ,int_R_DATA_TEMPR68[11] , 
       int_R_DATA_TEMPR68[10] ,int_R_DATA_TEMPR68[9] ,int_R_DATA_TEMPR68[8] , 
       int_R_DATA_TEMPR68[7] ,int_R_DATA_TEMPR68[6] ,int_R_DATA_TEMPR68[5] , 
       int_R_DATA_TEMPR68[4] ,int_R_DATA_TEMPR68[3] ,int_R_DATA_TEMPR68[2] , 
       int_R_DATA_TEMPR68[1] ,int_R_DATA_TEMPR68[0] }), .DB_DETECT( int_DB_DETECT_NG[68] ), .SB_CORRECT(int_SB_CORRECT_NG[68] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[68] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[17] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[17] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_16 (.A(sel_R_DATA_TEMPR16[31] ), .B(sel_R_DATA_TEMPR17[31] ), .C(sel_R_DATA_TEMPR18[31] ), .D(sel_R_DATA_TEMPR19[31] ), .Y(OR4_16_Y));
    OR4 OR4_386 (.A(sel_R_DATA_TEMPR28[21] ), .B(sel_R_DATA_TEMPR29[21] ), 
        .C(sel_R_DATA_TEMPR30[21] ), .D(sel_R_DATA_TEMPR31[21] ), .Y(
        OR4_386_Y));
    OR4 OR4_1327 (.A(OR4_955_Y), .B(OR4_734_Y), .C(OR4_502_Y), .D(
        OR4_519_Y), .Y(OR4_1327_Y));
    OR4 OR4_447 (.A(OR4_988_Y), .B(OR4_77_Y), .C(OR4_660_Y), .D(
        OR4_1246_Y), .Y(OR4_447_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%65%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R65C0 (.A_DOUT({
        nc584, nc585, nc586, nc587, nc588,int_R_DATA_TEMPR65[31] , 
       int_R_DATA_TEMPR65[30] ,int_R_DATA_TEMPR65[29] , 
       int_R_DATA_TEMPR65[28] ,int_R_DATA_TEMPR65[27] , 
       int_R_DATA_TEMPR65[26] ,int_R_DATA_TEMPR65[25] , 
       int_R_DATA_TEMPR65[24] ,int_R_DATA_TEMPR65[23] , 
       int_R_DATA_TEMPR65[22] ,int_R_DATA_TEMPR65[21] , 
       int_R_DATA_TEMPR65[20] ,int_R_DATA_TEMPR65[19] , 
       int_R_DATA_TEMPR65[18] ,int_R_DATA_TEMPR65[17] }), .B_DOUT({nc589, 
        nc590, nc591,int_R_DATA_TEMPR65[16] ,int_R_DATA_TEMPR65[15] , 
       int_R_DATA_TEMPR65[14] ,int_R_DATA_TEMPR65[13] , 
       int_R_DATA_TEMPR65[12] ,int_R_DATA_TEMPR65[11] , 
       int_R_DATA_TEMPR65[10] ,int_R_DATA_TEMPR65[9] ,int_R_DATA_TEMPR65[8] , 
       int_R_DATA_TEMPR65[7] ,int_R_DATA_TEMPR65[6] ,int_R_DATA_TEMPR65[5] , 
       int_R_DATA_TEMPR65[4] ,int_R_DATA_TEMPR65[3] ,int_R_DATA_TEMPR65[2] , 
       int_R_DATA_TEMPR65[1] ,int_R_DATA_TEMPR65[0] }), .DB_DETECT( int_DB_DETECT_NG[65] ), .SB_CORRECT(int_SB_CORRECT_NG[65] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[65] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[16] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[16] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_259 (.A(sel_R_DATA_TEMPR56[22] ), .B(sel_R_DATA_TEMPR57[22] ), 
        .C(sel_R_DATA_TEMPR58[22] ), .D(sel_R_DATA_TEMPR59[22] ), .Y(
        OR4_259_Y));
    OR4 OR4_4 (.A(sel_R_DATA_TEMPR96[27] ), .B(sel_R_DATA_TEMPR97[27] ), .C(sel_R_DATA_TEMPR98[27] ), .D(sel_R_DATA_TEMPR99[27] ), .Y(OR4_4_Y));
    OR4 OR4_331 (.A(OR4_417_Y), .B(OR4_856_Y), .C(OR4_1231_Y), .D(
        OR4_467_Y), .Y(OR4_331_Y));
    OR4 OR4_1171 (.A(OR4_1095_Y), .B(OR4_933_Y), .C(OR4_614_Y), .D(
        OR4_487_Y), .Y(OR4_1171_Y));
    OR4 OR4_512 (.A(sel_R_DATA_TEMPR124[16] ), .B(sel_R_DATA_TEMPR125[16] ), 
        .C(sel_R_DATA_TEMPR126[16] ), .D(sel_R_DATA_TEMPR127[16] ), .Y(
        OR4_512_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[4]  (.D(\BLKY2[4] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[4] ));
    OR4 OR4_1207 (.A(sel_R_DATA_TEMPR0[3] ), .B(sel_R_DATA_TEMPR1[3] ), .C(sel_R_DATA_TEMPR2[3] ), .D(sel_R_DATA_TEMPR3[3] ), .Y(OR4_1207_Y));
    OR4 OR4_320 (.A(sel_R_DATA_TEMPR4[31] ), .B(sel_R_DATA_TEMPR5[31] ), .C(sel_R_DATA_TEMPR6[31] ), .D(sel_R_DATA_TEMPR7[31] ), .Y(OR4_320_Y));
    OR4 OR4_430 (.A(sel_R_DATA_TEMPR20[6] ), .B(sel_R_DATA_TEMPR21[6] ), .C(sel_R_DATA_TEMPR22[6] ), .D(sel_R_DATA_TEMPR23[6] ), .Y(OR4_430_Y));
    OR4 OR4_1265 (.A(sel_R_DATA_TEMPR100[13] ), .B(sel_R_DATA_TEMPR101[13] ), 
        .C(sel_R_DATA_TEMPR102[13] ), .D(sel_R_DATA_TEMPR103[13] ), .Y(
        OR4_1265_Y));
    OR4 \OR4_R_DATA[14]  (.A(OR4_1316_Y), .B(OR4_822_Y), .C(OR4_113_Y), 
        .D(OR4_720_Y), .Y(R_DATA[14]));
    OR4 OR4_595 (.A(sel_R_DATA_TEMPR92[1] ), .B(sel_R_DATA_TEMPR93[1] ), .C(sel_R_DATA_TEMPR94[1] ), .D(sel_R_DATA_TEMPR95[1] ), .Y(OR4_595_Y));
    OR4 OR4_245 (.A(sel_R_DATA_TEMPR52[29] ), .B(sel_R_DATA_TEMPR53[29] ), 
        .C(sel_R_DATA_TEMPR54[29] ), .D(sel_R_DATA_TEMPR55[29] ), .Y(
        OR4_245_Y));
    OR4 OR4_508 (.A(OR4_0_Y), .B(OR2_20_Y), .C(sel_R_DATA_TEMPR86[11] ), 
        .D(sel_R_DATA_TEMPR87[11] ), .Y(OR4_508_Y));
    OR4 OR4_1390 (.A(sel_R_DATA_TEMPR56[12] ), .B(sel_R_DATA_TEMPR57[12] ), 
        .C(sel_R_DATA_TEMPR58[12] ), .D(sel_R_DATA_TEMPR59[12] ), .Y(
        OR4_1390_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[1]  (.D(\BLKY2[1] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[1] ));
    OR4 OR4_50 (.A(sel_R_DATA_TEMPR92[17] ), .B(sel_R_DATA_TEMPR93[17] ), .C(sel_R_DATA_TEMPR94[17] ), .D(sel_R_DATA_TEMPR95[17] ), .Y(OR4_50_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%42%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R42C0 (.A_DOUT({
        nc592, nc593, nc594, nc595, nc596,int_R_DATA_TEMPR42[31] , 
       int_R_DATA_TEMPR42[30] ,int_R_DATA_TEMPR42[29] , 
       int_R_DATA_TEMPR42[28] ,int_R_DATA_TEMPR42[27] , 
       int_R_DATA_TEMPR42[26] ,int_R_DATA_TEMPR42[25] , 
       int_R_DATA_TEMPR42[24] ,int_R_DATA_TEMPR42[23] , 
       int_R_DATA_TEMPR42[22] ,int_R_DATA_TEMPR42[21] , 
       int_R_DATA_TEMPR42[20] ,int_R_DATA_TEMPR42[19] , 
       int_R_DATA_TEMPR42[18] ,int_R_DATA_TEMPR42[17] }), .B_DOUT({nc597, 
        nc598, nc599,int_R_DATA_TEMPR42[16] ,int_R_DATA_TEMPR42[15] , 
       int_R_DATA_TEMPR42[14] ,int_R_DATA_TEMPR42[13] , 
       int_R_DATA_TEMPR42[12] ,int_R_DATA_TEMPR42[11] , 
       int_R_DATA_TEMPR42[10] ,int_R_DATA_TEMPR42[9] ,int_R_DATA_TEMPR42[8] , 
       int_R_DATA_TEMPR42[7] ,int_R_DATA_TEMPR42[6] ,int_R_DATA_TEMPR42[5] , 
       int_R_DATA_TEMPR42[4] ,int_R_DATA_TEMPR42[3] ,int_R_DATA_TEMPR42[2] , 
       int_R_DATA_TEMPR42[1] ,int_R_DATA_TEMPR42[0] }), .DB_DETECT( int_DB_DETECT_NG[42] ), .SB_CORRECT(int_SB_CORRECT_NG[42] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[42] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[10] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[10] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_842 (.A(\SB_CORRECT[60] ), .B(\SB_CORRECT[61] ), .C(
        \SB_CORRECT[62] ), .D(\SB_CORRECT[63] ), .Y(OR4_842_Y));
    OR4 OR4_1304 (.A(sel_R_DATA_TEMPR56[10] ), .B(sel_R_DATA_TEMPR57[10] ), 
        .C(sel_R_DATA_TEMPR58[10] ), .D(sel_R_DATA_TEMPR59[10] ), .Y(
        OR4_1304_Y));
    OR4 OR4_859 (.A(sel_R_DATA_TEMPR72[12] ), .B(sel_R_DATA_TEMPR73[12] ), 
        .C(sel_R_DATA_TEMPR74[12] ), .D(sel_R_DATA_TEMPR75[12] ), .Y(
        OR4_859_Y));
    OR4 OR4_823 (.A(sel_R_DATA_TEMPR64[10] ), .B(sel_R_DATA_TEMPR65[10] ), 
        .C(sel_R_DATA_TEMPR66[10] ), .D(sel_R_DATA_TEMPR67[10] ), .Y(
        OR4_823_Y));
    OR4 OR4_514 (.A(sel_R_DATA_TEMPR20[10] ), .B(sel_R_DATA_TEMPR21[10] ), 
        .C(sel_R_DATA_TEMPR22[10] ), .D(sel_R_DATA_TEMPR23[10] ), .Y(
        OR4_514_Y));
    OR4 OR4_1336 (.A(\SB_CORRECT[20] ), .B(\SB_CORRECT[21] ), .C(
        \SB_CORRECT[22] ), .D(\SB_CORRECT[23] ), .Y(OR4_1336_Y));
    OR4 OR4_578 (.A(OR4_136_Y), .B(OR4_895_Y), .C(OR4_1371_Y), .D(
        OR4_838_Y), .Y(OR4_578_Y));
    OR4 OR4_693 (.A(OR4_46_Y), .B(OR4_464_Y), .C(OR4_440_Y), .D(
        OR4_1097_Y), .Y(OR4_693_Y));
    OR4 OR4_57 (.A(sel_R_DATA_TEMPR0[12] ), .B(sel_R_DATA_TEMPR1[12] ), .C(sel_R_DATA_TEMPR2[12] ), .D(sel_R_DATA_TEMPR3[12] ), .Y(OR4_57_Y));
    AND4 \AND4DB_DETECT[33]  (.A(sel_DB_DETECT_NG[33] ), .B(
        \BLKY2_pipe[8] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[33] ));
    AND4 \AND4SB_CORRECT[32]  (.A(sel_SB_CORRECT_NG[32] ), .B(
        \BLKY2_pipe[8] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[32] ));
    OR4 OR4_32 (.A(sel_R_DATA_TEMPR24[0] ), .B(sel_R_DATA_TEMPR25[0] ), .C(sel_R_DATA_TEMPR26[0] ), .D(sel_R_DATA_TEMPR27[0] ), .Y(OR4_32_Y));
    OR4 OR4_260 (.A(sel_R_DATA_TEMPR28[0] ), .B(sel_R_DATA_TEMPR29[0] ), .C(sel_R_DATA_TEMPR30[0] ), .D(sel_R_DATA_TEMPR31[0] ), .Y(OR4_260_Y));
    OR4 OR4_912 (.A(OR4_36_Y), .B(OR4_308_Y), .C(OR4_1232_Y), .D(
        OR4_557_Y), .Y(OR4_912_Y));
    OR4 OR4_567 (.A(OR4_836_Y), .B(OR4_1344_Y), .C(OR4_608_Y), .D(
        OR4_827_Y), .Y(OR4_567_Y));
    OR4 OR4_1057 (.A(sel_R_DATA_TEMPR76[8] ), .B(sel_R_DATA_TEMPR77[8] ), .C(sel_R_DATA_TEMPR78[8] ), .D(sel_R_DATA_TEMPR79[8] ), .Y(OR4_1057_Y));
    AND4 \AND4SB_CORRECT[98]  (.A(sel_SB_CORRECT_NG[98] ), .B(
        \BLKY2_pipe[24] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[98] ));
    OR4 OR4_1287 (.A(sel_R_DATA_TEMPR28[24] ), .B(sel_R_DATA_TEMPR29[24] ), 
        .C(sel_R_DATA_TEMPR30[24] ), .D(sel_R_DATA_TEMPR31[24] ), .Y(
        OR4_1287_Y));
    OR4 OR4_406 (.A(sel_R_DATA_TEMPR48[20] ), .B(sel_R_DATA_TEMPR49[20] ), 
        .C(sel_R_DATA_TEMPR50[20] ), .D(sel_R_DATA_TEMPR51[20] ), .Y(
        OR4_406_Y));
    OR4 OR4_1016 (.A(sel_R_DATA_TEMPR68[15] ), .B(sel_R_DATA_TEMPR69[15] ), 
        .C(sel_R_DATA_TEMPR70[15] ), .D(sel_R_DATA_TEMPR71[15] ), .Y(
        OR4_1016_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%70%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R70C0 (.A_DOUT({
        nc600, nc601, nc602, nc603, nc604,int_R_DATA_TEMPR70[31] , 
       int_R_DATA_TEMPR70[30] ,int_R_DATA_TEMPR70[29] , 
       int_R_DATA_TEMPR70[28] ,int_R_DATA_TEMPR70[27] , 
       int_R_DATA_TEMPR70[26] ,int_R_DATA_TEMPR70[25] , 
       int_R_DATA_TEMPR70[24] ,int_R_DATA_TEMPR70[23] , 
       int_R_DATA_TEMPR70[22] ,int_R_DATA_TEMPR70[21] , 
       int_R_DATA_TEMPR70[20] ,int_R_DATA_TEMPR70[19] , 
       int_R_DATA_TEMPR70[18] ,int_R_DATA_TEMPR70[17] }), .B_DOUT({nc605, 
        nc606, nc607,int_R_DATA_TEMPR70[16] ,int_R_DATA_TEMPR70[15] , 
       int_R_DATA_TEMPR70[14] ,int_R_DATA_TEMPR70[13] , 
       int_R_DATA_TEMPR70[12] ,int_R_DATA_TEMPR70[11] , 
       int_R_DATA_TEMPR70[10] ,int_R_DATA_TEMPR70[9] ,int_R_DATA_TEMPR70[8] , 
       int_R_DATA_TEMPR70[7] ,int_R_DATA_TEMPR70[6] ,int_R_DATA_TEMPR70[5] , 
       int_R_DATA_TEMPR70[4] ,int_R_DATA_TEMPR70[3] ,int_R_DATA_TEMPR70[2] , 
       int_R_DATA_TEMPR70[1] ,int_R_DATA_TEMPR70[0] }), .DB_DETECT( int_DB_DETECT_NG[70] ), .SB_CORRECT(int_SB_CORRECT_NG[70] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[70] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[17] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[17] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1075 (.A(\SB_CORRECT[72] ), .B(\SB_CORRECT[73] ), .C(
        \SB_CORRECT[74] ), .D(\SB_CORRECT[75] ), .Y(OR4_1075_Y));
    OR4 OR4_443 (.A(sel_R_DATA_TEMPR112[6] ), .B(sel_R_DATA_TEMPR113[6] ), 
        .C(sel_R_DATA_TEMPR114[6] ), .D(sel_R_DATA_TEMPR115[6] ), .Y(
        OR4_443_Y));
    OR4 OR4_669 (.A(sel_R_DATA_TEMPR16[10] ), .B(sel_R_DATA_TEMPR17[10] ), 
        .C(sel_R_DATA_TEMPR18[10] ), .D(sel_R_DATA_TEMPR19[10] ), .Y(
        OR4_669_Y));
    OR4 OR4_641 (.A(sel_R_DATA_TEMPR48[18] ), .B(sel_R_DATA_TEMPR49[18] ), 
        .C(sel_R_DATA_TEMPR50[18] ), .D(sel_R_DATA_TEMPR51[18] ), .Y(
        OR4_641_Y));
    OR4 OR4_476 (.A(sel_R_DATA_TEMPR60[22] ), .B(sel_R_DATA_TEMPR61[22] ), 
        .C(sel_R_DATA_TEMPR62[22] ), .D(sel_R_DATA_TEMPR63[22] ), .Y(
        OR4_476_Y));
    OR4 OR4_184 (.A(sel_R_DATA_TEMPR20[25] ), .B(sel_R_DATA_TEMPR21[25] ), 
        .C(sel_R_DATA_TEMPR22[25] ), .D(sel_R_DATA_TEMPR23[25] ), .Y(
        OR4_184_Y));
    OR4 OR4_311 (.A(sel_R_DATA_TEMPR60[0] ), .B(sel_R_DATA_TEMPR61[0] ), .C(sel_R_DATA_TEMPR62[0] ), .D(sel_R_DATA_TEMPR63[0] ), .Y(OR4_311_Y));
    AND4 \AND4SB_CORRECT[110]  (.A(sel_SB_CORRECT_NG[110] ), .B(
        \BLKY2_pipe[27] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[110] ));
    AND4 \AND4SB_CORRECT[15]  (.A(sel_SB_CORRECT_NG[15] ), .B(
        \BLKY2_pipe[3] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[15] ));
    AND4 \AND4SB_CORRECT[16]  (.A(sel_SB_CORRECT_NG[16] ), .B(
        \BLKY2_pipe[4] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[16] ));
    OR4 OR4_248 (.A(sel_R_DATA_TEMPR108[7] ), .B(sel_R_DATA_TEMPR109[7] ), 
        .C(sel_R_DATA_TEMPR110[7] ), .D(sel_R_DATA_TEMPR111[7] ), .Y(
        OR4_248_Y));
    OR4 OR4_1384 (.A(sel_R_DATA_TEMPR72[5] ), .B(sel_R_DATA_TEMPR73[5] ), .C(sel_R_DATA_TEMPR74[5] ), .D(sel_R_DATA_TEMPR75[5] ), .Y(OR4_1384_Y));
    OR4 OR4_999 (.A(sel_R_DATA_TEMPR108[9] ), .B(sel_R_DATA_TEMPR109[9] ), 
        .C(sel_R_DATA_TEMPR110[9] ), .D(sel_R_DATA_TEMPR111[9] ), .Y(
        OR4_999_Y));
    OR4 OR4_990 (.A(OR4_416_Y), .B(OR4_891_Y), .C(OR4_1366_Y), .D(
        OR4_354_Y), .Y(OR4_990_Y));
    OR4 OR4_1311 (.A(OR4_448_Y), .B(OR4_691_Y), .C(OR4_900_Y), .D(
        OR4_739_Y), .Y(OR4_1311_Y));
    OR4 OR4_757 (.A(OR4_639_Y), .B(OR2_2_Y), .C(sel_R_DATA_TEMPR86[25] ), 
        .D(sel_R_DATA_TEMPR87[25] ), .Y(OR4_757_Y));
    OR4 OR4_1309 (.A(sel_R_DATA_TEMPR104[29] ), .B(sel_R_DATA_TEMPR105[29] ), 
        .C(sel_R_DATA_TEMPR106[29] ), .D(sel_R_DATA_TEMPR107[29] ), .Y(
        OR4_1309_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%1%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R1C0 (.A_DOUT({
        nc608, nc609, nc610, nc611, nc612,int_R_DATA_TEMPR1[31] , 
       int_R_DATA_TEMPR1[30] ,int_R_DATA_TEMPR1[29] ,int_R_DATA_TEMPR1[28] , 
       int_R_DATA_TEMPR1[27] ,int_R_DATA_TEMPR1[26] ,int_R_DATA_TEMPR1[25] , 
       int_R_DATA_TEMPR1[24] ,int_R_DATA_TEMPR1[23] ,int_R_DATA_TEMPR1[22] , 
       int_R_DATA_TEMPR1[21] ,int_R_DATA_TEMPR1[20] ,int_R_DATA_TEMPR1[19] , 
       int_R_DATA_TEMPR1[18] ,int_R_DATA_TEMPR1[17] }), .B_DOUT({nc613, 
        nc614, nc615,int_R_DATA_TEMPR1[16] ,int_R_DATA_TEMPR1[15] , 
       int_R_DATA_TEMPR1[14] ,int_R_DATA_TEMPR1[13] ,int_R_DATA_TEMPR1[12] , 
       int_R_DATA_TEMPR1[11] ,int_R_DATA_TEMPR1[10] ,int_R_DATA_TEMPR1[9] , 
       int_R_DATA_TEMPR1[8] ,int_R_DATA_TEMPR1[7] ,int_R_DATA_TEMPR1[6] , 
       int_R_DATA_TEMPR1[5] ,int_R_DATA_TEMPR1[4] ,int_R_DATA_TEMPR1[3] , 
       int_R_DATA_TEMPR1[2] ,int_R_DATA_TEMPR1[1] ,int_R_DATA_TEMPR1[0] }), 
        .DB_DETECT(int_DB_DETECT_NG[1] ), .SB_CORRECT( int_SB_CORRECT_NG[1] ), .ACCESS_BUSY(\ACCESS_BUSY[1] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[0] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[30]  (.A(CFG3_1_Y), .B(CFG3_3_Y)
        , .Y(\BLKY2[30] ));
    OR4 OR4_754 (.A(sel_R_DATA_TEMPR32[4] ), .B(sel_R_DATA_TEMPR33[4] ), .C(sel_R_DATA_TEMPR34[4] ), .D(sel_R_DATA_TEMPR35[4] ), .Y(OR4_754_Y));
    OR4 OR4_302 (.A(sel_R_DATA_TEMPR116[17] ), .B(sel_R_DATA_TEMPR117[17] ), 
        .C(sel_R_DATA_TEMPR118[17] ), .D(sel_R_DATA_TEMPR119[17] ), .Y(
        OR4_302_Y));
    OR4 OR4_266 (.A(OR4_780_Y), .B(OR4_1053_Y), .C(OR4_1269_Y), .D(
        OR4_1098_Y), .Y(OR4_266_Y));
    OR4 OR4_SB_CORRECT (.A(OR4_518_Y), .B(OR4_1263_Y), .C(OR4_765_Y), 
        .D(OR4_256_Y), .Y(SB_CORRECT));
    AND4 \AND4DB_DETECT[15]  (.A(sel_DB_DETECT_NG[15] ), .B(
        \BLKY2_pipe[3] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[15] ));
    OR4 OR4_1295 (.A(\DB_DETECT[24] ), .B(\DB_DETECT[25] ), .C(
        \DB_DETECT[26] ), .D(\DB_DETECT[27] ), .Y(OR4_1295_Y));
    AND4 \AND4SB_CORRECT[73]  (.A(sel_SB_CORRECT_NG[73] ), .B(
        \BLKY2_pipe[18] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[73] ));
    OR4 OR4_1000 (.A(sel_R_DATA_TEMPR52[4] ), .B(sel_R_DATA_TEMPR53[4] ), .C(sel_R_DATA_TEMPR54[4] ), .D(sel_R_DATA_TEMPR55[4] ), .Y(OR4_1000_Y));
    OR4 OR4_10 (.A(sel_R_DATA_TEMPR40[1] ), .B(sel_R_DATA_TEMPR41[1] ), .C(sel_R_DATA_TEMPR42[1] ), .D(sel_R_DATA_TEMPR43[1] ), .Y(OR4_10_Y));
    OR4 OR4_25 (.A(sel_R_DATA_TEMPR100[12] ), .B(sel_R_DATA_TEMPR101[12] ), 
        .C(sel_R_DATA_TEMPR102[12] ), .D(sel_R_DATA_TEMPR103[12] ), .Y(
        OR4_25_Y));
    OR4 OR4_76 (.A(sel_R_DATA_TEMPR80[27] ), .B(sel_R_DATA_TEMPR81[27] ), .C(sel_R_DATA_TEMPR82[27] ), .D(sel_R_DATA_TEMPR83[27] ), .Y(OR4_76_Y));
    OR4 OR4_410 (.A(OR4_405_Y), .B(OR2_30_Y), .C(sel_R_DATA_TEMPR86[23] ), 
        .D(sel_R_DATA_TEMPR87[23] ), .Y(OR4_410_Y));
    OR4 OR4_983 (.A(sel_R_DATA_TEMPR56[24] ), .B(sel_R_DATA_TEMPR57[24] ), 
        .C(sel_R_DATA_TEMPR58[24] ), .D(sel_R_DATA_TEMPR59[24] ), .Y(
        OR4_983_Y));
    OR4 OR4_339 (.A(sel_R_DATA_TEMPR4[8] ), .B(sel_R_DATA_TEMPR5[8] ), .C(sel_R_DATA_TEMPR6[8] ), .D(sel_R_DATA_TEMPR7[8] ), .Y(OR4_339_Y));
    OR4 OR4_193 (.A(sel_R_DATA_TEMPR44[20] ), .B(sel_R_DATA_TEMPR45[20] ), 
        .C(sel_R_DATA_TEMPR46[20] ), .D(sel_R_DATA_TEMPR47[20] ), .Y(
        OR4_193_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%14%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R14C0 (.A_DOUT({
        nc616, nc617, nc618, nc619, nc620,int_R_DATA_TEMPR14[31] , 
       int_R_DATA_TEMPR14[30] ,int_R_DATA_TEMPR14[29] , 
       int_R_DATA_TEMPR14[28] ,int_R_DATA_TEMPR14[27] , 
       int_R_DATA_TEMPR14[26] ,int_R_DATA_TEMPR14[25] , 
       int_R_DATA_TEMPR14[24] ,int_R_DATA_TEMPR14[23] , 
       int_R_DATA_TEMPR14[22] ,int_R_DATA_TEMPR14[21] , 
       int_R_DATA_TEMPR14[20] ,int_R_DATA_TEMPR14[19] , 
       int_R_DATA_TEMPR14[18] ,int_R_DATA_TEMPR14[17] }), .B_DOUT({nc621, 
        nc622, nc623,int_R_DATA_TEMPR14[16] ,int_R_DATA_TEMPR14[15] , 
       int_R_DATA_TEMPR14[14] ,int_R_DATA_TEMPR14[13] , 
       int_R_DATA_TEMPR14[12] ,int_R_DATA_TEMPR14[11] , 
       int_R_DATA_TEMPR14[10] ,int_R_DATA_TEMPR14[9] ,int_R_DATA_TEMPR14[8] , 
       int_R_DATA_TEMPR14[7] ,int_R_DATA_TEMPR14[6] ,int_R_DATA_TEMPR14[5] , 
       int_R_DATA_TEMPR14[4] ,int_R_DATA_TEMPR14[3] ,int_R_DATA_TEMPR14[2] , 
       int_R_DATA_TEMPR14[1] ,int_R_DATA_TEMPR14[0] }), .DB_DETECT( int_DB_DETECT_NG[14] ), .SB_CORRECT(int_SB_CORRECT_NG[14] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[14] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[3] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_372 (.A(OR4_901_Y), .B(OR4_761_Y), .C(OR4_859_Y), .D(
        OR4_644_Y), .Y(OR4_372_Y));
    OR4 OR4_1246 (.A(OR4_187_Y), .B(OR4_460_Y), .C(OR4_648_Y), .D(
        OR4_497_Y), .Y(OR4_1246_Y));
    OR4 OR4_851 (.A(sel_R_DATA_TEMPR88[23] ), .B(sel_R_DATA_TEMPR89[23] ), 
        .C(sel_R_DATA_TEMPR90[23] ), .D(sel_R_DATA_TEMPR91[23] ), .Y(
        OR4_851_Y));
    OR4 OR4_525 (.A(OR4_1208_Y), .B(OR4_773_Y), .C(OR4_848_Y), .D(
        OR4_1111_Y), .Y(OR4_525_Y));
    OR4 OR4_17 (.A(OR4_5_Y), .B(OR4_725_Y), .C(OR4_18_Y), .D(OR4_241_Y)
        , .Y(OR4_17_Y));
    OR4 OR4_886 (.A(sel_R_DATA_TEMPR100[3] ), .B(sel_R_DATA_TEMPR101[3] ), 
        .C(sel_R_DATA_TEMPR102[3] ), .D(sel_R_DATA_TEMPR103[3] ), .Y(
        OR4_886_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%81%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R81C0 (.A_DOUT({
        nc624, nc625, nc626, nc627, nc628,int_R_DATA_TEMPR81[31] , 
       int_R_DATA_TEMPR81[30] ,int_R_DATA_TEMPR81[29] , 
       int_R_DATA_TEMPR81[28] ,int_R_DATA_TEMPR81[27] , 
       int_R_DATA_TEMPR81[26] ,int_R_DATA_TEMPR81[25] , 
       int_R_DATA_TEMPR81[24] ,int_R_DATA_TEMPR81[23] , 
       int_R_DATA_TEMPR81[22] ,int_R_DATA_TEMPR81[21] , 
       int_R_DATA_TEMPR81[20] ,int_R_DATA_TEMPR81[19] , 
       int_R_DATA_TEMPR81[18] ,int_R_DATA_TEMPR81[17] }), .B_DOUT({nc629, 
        nc630, nc631,int_R_DATA_TEMPR81[16] ,int_R_DATA_TEMPR81[15] , 
       int_R_DATA_TEMPR81[14] ,int_R_DATA_TEMPR81[13] , 
       int_R_DATA_TEMPR81[12] ,int_R_DATA_TEMPR81[11] , 
       int_R_DATA_TEMPR81[10] ,int_R_DATA_TEMPR81[9] ,int_R_DATA_TEMPR81[8] , 
       int_R_DATA_TEMPR81[7] ,int_R_DATA_TEMPR81[6] ,int_R_DATA_TEMPR81[5] , 
       int_R_DATA_TEMPR81[4] ,int_R_DATA_TEMPR81[3] ,int_R_DATA_TEMPR81[2] , 
       int_R_DATA_TEMPR81[1] ,int_R_DATA_TEMPR81[0] }), .DB_DETECT( int_DB_DETECT_NG[81] ), .SB_CORRECT(int_SB_CORRECT_NG[81] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[81] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[20] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[20] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_781 (.A(OR4_524_Y), .B(OR2_28_Y), .C(sel_R_DATA_TEMPR86[17] ), 
        .D(sel_R_DATA_TEMPR87[17] ), .Y(OR4_781_Y));
    OR4 OR4_664 (.A(\DB_DETECT[4] ), .B(\DB_DETECT[5] ), .C(
        \DB_DETECT[6] ), .D(\DB_DETECT[7] ), .Y(OR4_664_Y));
    OR4 OR4_1326 (.A(sel_R_DATA_TEMPR88[13] ), .B(sel_R_DATA_TEMPR89[13] ), 
        .C(sel_R_DATA_TEMPR90[13] ), .D(sel_R_DATA_TEMPR91[13] ), .Y(
        OR4_1326_Y));
    OR4 OR4_1348 (.A(sel_R_DATA_TEMPR0[8] ), .B(sel_R_DATA_TEMPR1[8] ), .C(sel_R_DATA_TEMPR2[8] ), .D(sel_R_DATA_TEMPR3[8] ), .Y(OR4_1348_Y));
    CFG3 #( .INIT(8'h4) )  CFG3_14 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_14_Y));
    OR4 OR4_623 (.A(sel_R_DATA_TEMPR8[15] ), .B(sel_R_DATA_TEMPR9[15] ), .C(sel_R_DATA_TEMPR10[15] ), .D(sel_R_DATA_TEMPR11[15] ), .Y(OR4_623_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%104%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R104C0 (.A_DOUT({
        nc632, nc633, nc634, nc635, nc636,int_R_DATA_TEMPR104[31] , 
       int_R_DATA_TEMPR104[30] ,int_R_DATA_TEMPR104[29] , 
       int_R_DATA_TEMPR104[28] ,int_R_DATA_TEMPR104[27] , 
       int_R_DATA_TEMPR104[26] ,int_R_DATA_TEMPR104[25] , 
       int_R_DATA_TEMPR104[24] ,int_R_DATA_TEMPR104[23] , 
       int_R_DATA_TEMPR104[22] ,int_R_DATA_TEMPR104[21] , 
       int_R_DATA_TEMPR104[20] ,int_R_DATA_TEMPR104[19] , 
       int_R_DATA_TEMPR104[18] ,int_R_DATA_TEMPR104[17] }), .B_DOUT({nc637, 
        nc638, nc639,int_R_DATA_TEMPR104[16] ,int_R_DATA_TEMPR104[15] , 
       int_R_DATA_TEMPR104[14] ,int_R_DATA_TEMPR104[13] , 
       int_R_DATA_TEMPR104[12] ,int_R_DATA_TEMPR104[11] , 
       int_R_DATA_TEMPR104[10] ,int_R_DATA_TEMPR104[9] , 
       int_R_DATA_TEMPR104[8] ,int_R_DATA_TEMPR104[7] , 
       int_R_DATA_TEMPR104[6] ,int_R_DATA_TEMPR104[5] , 
       int_R_DATA_TEMPR104[4] ,int_R_DATA_TEMPR104[3] , 
       int_R_DATA_TEMPR104[2] ,int_R_DATA_TEMPR104[1] , 
       int_R_DATA_TEMPR104[0] }), .DB_DETECT(int_DB_DETECT_NG[104] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[104] ), .ACCESS_BUSY(
        ACCESS_BUSY[104] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[26] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[26] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1389 (.A(sel_R_DATA_TEMPR108[27] ), .B(sel_R_DATA_TEMPR109[27] ), 
        .C(sel_R_DATA_TEMPR110[27] ), .D(sel_R_DATA_TEMPR111[27] ), .Y(
        OR4_1389_Y));
    AND4 \AND4DB_DETECT[96]  (.A(sel_DB_DETECT_NG[96] ), .B(
        \BLKY2_pipe[24] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[96] ));
    AND4 \AND4SB_CORRECT[74]  (.A(sel_SB_CORRECT_NG[74] ), .B(
        \BLKY2_pipe[18] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[74] ));
    OR4 OR4_586 (.A(OR4_55_Y), .B(OR4_1291_Y), .C(OR4_767_Y), .D(
        OR4_1234_Y), .Y(OR4_586_Y));
    OR4 OR4_1080 (.A(OR4_1268_Y), .B(OR4_1147_Y), .C(OR4_1075_Y), .D(
        OR4_663_Y), .Y(OR4_1080_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%32%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R32C0 (.A_DOUT({
        nc640, nc641, nc642, nc643, nc644,int_R_DATA_TEMPR32[31] , 
       int_R_DATA_TEMPR32[30] ,int_R_DATA_TEMPR32[29] , 
       int_R_DATA_TEMPR32[28] ,int_R_DATA_TEMPR32[27] , 
       int_R_DATA_TEMPR32[26] ,int_R_DATA_TEMPR32[25] , 
       int_R_DATA_TEMPR32[24] ,int_R_DATA_TEMPR32[23] , 
       int_R_DATA_TEMPR32[22] ,int_R_DATA_TEMPR32[21] , 
       int_R_DATA_TEMPR32[20] ,int_R_DATA_TEMPR32[19] , 
       int_R_DATA_TEMPR32[18] ,int_R_DATA_TEMPR32[17] }), .B_DOUT({nc645, 
        nc646, nc647,int_R_DATA_TEMPR32[16] ,int_R_DATA_TEMPR32[15] , 
       int_R_DATA_TEMPR32[14] ,int_R_DATA_TEMPR32[13] , 
       int_R_DATA_TEMPR32[12] ,int_R_DATA_TEMPR32[11] , 
       int_R_DATA_TEMPR32[10] ,int_R_DATA_TEMPR32[9] ,int_R_DATA_TEMPR32[8] , 
       int_R_DATA_TEMPR32[7] ,int_R_DATA_TEMPR32[6] ,int_R_DATA_TEMPR32[5] , 
       int_R_DATA_TEMPR32[4] ,int_R_DATA_TEMPR32[3] ,int_R_DATA_TEMPR32[2] , 
       int_R_DATA_TEMPR32[1] ,int_R_DATA_TEMPR32[0] }), .DB_DETECT( int_DB_DETECT_NG[32] ), .SB_CORRECT(int_SB_CORRECT_NG[32] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[32] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[8] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[8] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1134 (.A(sel_R_DATA_TEMPR4[4] ), .B(sel_R_DATA_TEMPR5[4] ), .C(sel_R_DATA_TEMPR6[4] ), .D(sel_R_DATA_TEMPR7[4] ), .Y(OR4_1134_Y));
    DFN1E1 \DFN1E1BLKY0_pipe[1]  (.D(R_ADDR[9]), .CLK(CLK), .E(VCC), 
        .Q(\BLKY0_pipe[1] ));
    AND4 \AND4DB_DETECT[91]  (.A(sel_DB_DETECT_NG[91] ), .B(
        \BLKY2_pipe[22] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[91] ));
    AND4 \AND4SB_CORRECT[80]  (.A(sel_SB_CORRECT_NG[80] ), .B(
        \BLKY2_pipe[20] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[80] ));
    DFN1E1 \DFN1E1BLKY2_pipe[7]  (.D(\BLKY2[7] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[7] ));
    OR4 OR4_200 (.A(sel_R_DATA_TEMPR108[10] ), .B(sel_R_DATA_TEMPR109[10] ), 
        .C(sel_R_DATA_TEMPR110[10] ), .D(sel_R_DATA_TEMPR111[10] ), .Y(
        OR4_200_Y));
    OR4 OR4_1064 (.A(sel_R_DATA_TEMPR92[14] ), .B(sel_R_DATA_TEMPR93[14] ), 
        .C(sel_R_DATA_TEMPR94[14] ), .D(sel_R_DATA_TEMPR95[14] ), .Y(
        OR4_1064_Y));
    OR4 OR4_507 (.A(sel_R_DATA_TEMPR56[25] ), .B(sel_R_DATA_TEMPR57[25] ), 
        .C(sel_R_DATA_TEMPR58[25] ), .D(sel_R_DATA_TEMPR59[25] ), .Y(
        OR4_507_Y));
    AND4 \AND4DB_DETECT[54]  (.A(sel_DB_DETECT_NG[54] ), .B(
        \BLKY2_pipe[13] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[54] ));
    AND4 \AND4DB_DETECT[66]  (.A(sel_DB_DETECT_NG[66] ), .B(
        \BLKY2_pipe[16] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[66] ));
    OR4 OR4_1049 (.A(sel_R_DATA_TEMPR120[23] ), .B(sel_R_DATA_TEMPR121[23] ), 
        .C(sel_R_DATA_TEMPR122[23] ), .D(sel_R_DATA_TEMPR123[23] ), .Y(
        OR4_1049_Y));
    OR4 OR4_270 (.A(sel_R_DATA_TEMPR12[20] ), .B(sel_R_DATA_TEMPR13[20] ), 
        .C(sel_R_DATA_TEMPR14[20] ), .D(sel_R_DATA_TEMPR15[20] ), .Y(
        OR4_270_Y));
    OR4 OR4_1363 (.A(OR4_1187_Y), .B(OR4_1374_Y), .C(OR4_1357_Y), .D(
        OR4_1072_Y), .Y(OR4_1363_Y));
    OR4 OR4_1170 (.A(sel_R_DATA_TEMPR12[22] ), .B(sel_R_DATA_TEMPR13[22] ), 
        .C(sel_R_DATA_TEMPR14[22] ), .D(sel_R_DATA_TEMPR15[22] ), .Y(
        OR4_1170_Y));
    OR4 OR4_929 (.A(OR4_103_Y), .B(OR4_370_Y), .C(OR4_566_Y), .D(
        OR4_414_Y), .Y(OR4_929_Y));
    OR4 OR4_920 (.A(sel_R_DATA_TEMPR112[7] ), .B(sel_R_DATA_TEMPR113[7] ), 
        .C(sel_R_DATA_TEMPR114[7] ), .D(sel_R_DATA_TEMPR115[7] ), .Y(
        OR4_920_Y));
    AND4 \AND4DB_DETECT[61]  (.A(sel_DB_DETECT_NG[61] ), .B(
        \BLKY2_pipe[15] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[61] ));
    OR4 OR4_890 (.A(sel_R_DATA_TEMPR72[20] ), .B(sel_R_DATA_TEMPR73[20] ), 
        .C(sel_R_DATA_TEMPR74[20] ), .D(sel_R_DATA_TEMPR75[20] ), .Y(
        OR4_890_Y));
    AND4 \AND4SB_CORRECT[53]  (.A(sel_SB_CORRECT_NG[53] ), .B(
        \BLKY2_pipe[13] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[53] ));
    OR4 OR4_577 (.A(OR4_784_Y), .B(OR4_375_Y), .C(OR4_425_Y), .D(
        OR4_824_Y), .Y(OR4_577_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[12]  (.A(CFG3_18_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[12] ));
    OR4 OR4_957 (.A(\DB_DETECT[88] ), .B(\DB_DETECT[89] ), .C(
        \DB_DETECT[90] ), .D(\DB_DETECT[91] ), .Y(OR4_957_Y));
    AND4 \AND4SB_CORRECT[49]  (.A(sel_SB_CORRECT_NG[49] ), .B(
        \BLKY2_pipe[12] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[49] ));
    OR4 OR4_739 (.A(sel_R_DATA_TEMPR108[17] ), .B(sel_R_DATA_TEMPR109[17] ), 
        .C(sel_R_DATA_TEMPR110[17] ), .D(sel_R_DATA_TEMPR111[17] ), .Y(
        OR4_739_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[21]  (.A(CFG3_22_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[21] ));
    OR4 OR4_541 (.A(sel_R_DATA_TEMPR36[8] ), .B(sel_R_DATA_TEMPR37[8] ), .C(sel_R_DATA_TEMPR38[8] ), .D(sel_R_DATA_TEMPR39[8] ), .Y(OR4_541_Y));
    OR4 OR4_192 (.A(sel_R_DATA_TEMPR108[2] ), .B(sel_R_DATA_TEMPR109[2] ), 
        .C(sel_R_DATA_TEMPR110[2] ), .D(sel_R_DATA_TEMPR111[2] ), .Y(
        OR4_192_Y));
    OR4 OR4_319 (.A(OR4_1105_Y), .B(OR2_9_Y), .C(sel_R_DATA_TEMPR86[15] ), 
        .D(sel_R_DATA_TEMPR87[15] ), .Y(OR4_319_Y));
    OR4 OR4_1238 (.A(sel_R_DATA_TEMPR48[24] ), .B(sel_R_DATA_TEMPR49[24] ), 
        .C(sel_R_DATA_TEMPR50[24] ), .D(sel_R_DATA_TEMPR51[24] ), .Y(
        OR4_1238_Y));
    OR4 OR4_609 (.A(sel_R_DATA_TEMPR16[28] ), .B(sel_R_DATA_TEMPR17[28] ), 
        .C(sel_R_DATA_TEMPR18[28] ), .D(sel_R_DATA_TEMPR19[28] ), .Y(
        OR4_609_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%27%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R27C0 (.A_DOUT({
        nc648, nc649, nc650, nc651, nc652,int_R_DATA_TEMPR27[31] , 
       int_R_DATA_TEMPR27[30] ,int_R_DATA_TEMPR27[29] , 
       int_R_DATA_TEMPR27[28] ,int_R_DATA_TEMPR27[27] , 
       int_R_DATA_TEMPR27[26] ,int_R_DATA_TEMPR27[25] , 
       int_R_DATA_TEMPR27[24] ,int_R_DATA_TEMPR27[23] , 
       int_R_DATA_TEMPR27[22] ,int_R_DATA_TEMPR27[21] , 
       int_R_DATA_TEMPR27[20] ,int_R_DATA_TEMPR27[19] , 
       int_R_DATA_TEMPR27[18] ,int_R_DATA_TEMPR27[17] }), .B_DOUT({nc653, 
        nc654, nc655,int_R_DATA_TEMPR27[16] ,int_R_DATA_TEMPR27[15] , 
       int_R_DATA_TEMPR27[14] ,int_R_DATA_TEMPR27[13] , 
       int_R_DATA_TEMPR27[12] ,int_R_DATA_TEMPR27[11] , 
       int_R_DATA_TEMPR27[10] ,int_R_DATA_TEMPR27[9] ,int_R_DATA_TEMPR27[8] , 
       int_R_DATA_TEMPR27[7] ,int_R_DATA_TEMPR27[6] ,int_R_DATA_TEMPR27[5] , 
       int_R_DATA_TEMPR27[4] ,int_R_DATA_TEMPR27[3] ,int_R_DATA_TEMPR27[2] , 
       int_R_DATA_TEMPR27[1] ,int_R_DATA_TEMPR27[0] }), .DB_DETECT( int_DB_DETECT_NG[27] ), .SB_CORRECT(int_SB_CORRECT_NG[27] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[27] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[6] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_995 (.A(sel_R_DATA_TEMPR12[9] ), .B(sel_R_DATA_TEMPR13[9] ), .C(sel_R_DATA_TEMPR14[9] ), .D(sel_R_DATA_TEMPR15[9] ), .Y(OR4_995_Y));
    OR4 OR4_123 (.A(sel_R_DATA_TEMPR72[27] ), .B(sel_R_DATA_TEMPR73[27] ), 
        .C(sel_R_DATA_TEMPR74[27] ), .D(sel_R_DATA_TEMPR75[27] ), .Y(
        OR4_123_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%58%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R58C0 (.A_DOUT({
        nc656, nc657, nc658, nc659, nc660,int_R_DATA_TEMPR58[31] , 
       int_R_DATA_TEMPR58[30] ,int_R_DATA_TEMPR58[29] , 
       int_R_DATA_TEMPR58[28] ,int_R_DATA_TEMPR58[27] , 
       int_R_DATA_TEMPR58[26] ,int_R_DATA_TEMPR58[25] , 
       int_R_DATA_TEMPR58[24] ,int_R_DATA_TEMPR58[23] , 
       int_R_DATA_TEMPR58[22] ,int_R_DATA_TEMPR58[21] , 
       int_R_DATA_TEMPR58[20] ,int_R_DATA_TEMPR58[19] , 
       int_R_DATA_TEMPR58[18] ,int_R_DATA_TEMPR58[17] }), .B_DOUT({nc661, 
        nc662, nc663,int_R_DATA_TEMPR58[16] ,int_R_DATA_TEMPR58[15] , 
       int_R_DATA_TEMPR58[14] ,int_R_DATA_TEMPR58[13] , 
       int_R_DATA_TEMPR58[12] ,int_R_DATA_TEMPR58[11] , 
       int_R_DATA_TEMPR58[10] ,int_R_DATA_TEMPR58[9] ,int_R_DATA_TEMPR58[8] , 
       int_R_DATA_TEMPR58[7] ,int_R_DATA_TEMPR58[6] ,int_R_DATA_TEMPR58[5] , 
       int_R_DATA_TEMPR58[4] ,int_R_DATA_TEMPR58[3] ,int_R_DATA_TEMPR58[2] , 
       int_R_DATA_TEMPR58[1] ,int_R_DATA_TEMPR58[0] }), .DB_DETECT( int_DB_DETECT_NG[58] ), .SB_CORRECT(int_SB_CORRECT_NG[58] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[58] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[14] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[14] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_834 (.A(OR4_265_Y), .B(OR4_559_Y), .C(OR4_1015_Y), .D(
        OR4_509_Y), .Y(OR4_834_Y));
    OR4 OR4_679 (.A(OR4_922_Y), .B(OR4_772_Y), .C(OR4_1252_Y), .D(
        OR4_239_Y), .Y(OR4_679_Y));
    OR4 OR4_1257 (.A(sel_R_DATA_TEMPR32[18] ), .B(sel_R_DATA_TEMPR33[18] ), 
        .C(sel_R_DATA_TEMPR34[18] ), .D(sel_R_DATA_TEMPR35[18] ), .Y(
        OR4_1257_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[2]  (.A(CFG3_14_Y), .B(
        CFG3_12_Y), .Y(\BLKX2[2] ));
    OR4 OR4_206 (.A(OR4_1174_Y), .B(OR4_857_Y), .C(OR4_1334_Y), .D(
        OR4_805_Y), .Y(OR4_206_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%55%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R55C0 (.A_DOUT({
        nc664, nc665, nc666, nc667, nc668,int_R_DATA_TEMPR55[31] , 
       int_R_DATA_TEMPR55[30] ,int_R_DATA_TEMPR55[29] , 
       int_R_DATA_TEMPR55[28] ,int_R_DATA_TEMPR55[27] , 
       int_R_DATA_TEMPR55[26] ,int_R_DATA_TEMPR55[25] , 
       int_R_DATA_TEMPR55[24] ,int_R_DATA_TEMPR55[23] , 
       int_R_DATA_TEMPR55[22] ,int_R_DATA_TEMPR55[21] , 
       int_R_DATA_TEMPR55[20] ,int_R_DATA_TEMPR55[19] , 
       int_R_DATA_TEMPR55[18] ,int_R_DATA_TEMPR55[17] }), .B_DOUT({nc669, 
        nc670, nc671,int_R_DATA_TEMPR55[16] ,int_R_DATA_TEMPR55[15] , 
       int_R_DATA_TEMPR55[14] ,int_R_DATA_TEMPR55[13] , 
       int_R_DATA_TEMPR55[12] ,int_R_DATA_TEMPR55[11] , 
       int_R_DATA_TEMPR55[10] ,int_R_DATA_TEMPR55[9] ,int_R_DATA_TEMPR55[8] , 
       int_R_DATA_TEMPR55[7] ,int_R_DATA_TEMPR55[6] ,int_R_DATA_TEMPR55[5] , 
       int_R_DATA_TEMPR55[4] ,int_R_DATA_TEMPR55[3] ,int_R_DATA_TEMPR55[2] , 
       int_R_DATA_TEMPR55[1] ,int_R_DATA_TEMPR55[0] }), .DB_DETECT( int_DB_DETECT_NG[55] ), .SB_CORRECT(int_SB_CORRECT_NG[55] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[55] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[13] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[13] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_533 (.A(sel_R_DATA_TEMPR0[10] ), .B(sel_R_DATA_TEMPR1[10] ), .C(sel_R_DATA_TEMPR2[10] ), .D(sel_R_DATA_TEMPR3[10] ), .Y(OR4_533_Y));
    OR4 OR4_70 (.A(sel_R_DATA_TEMPR64[31] ), .B(sel_R_DATA_TEMPR65[31] ), .C(sel_R_DATA_TEMPR66[31] ), .D(sel_R_DATA_TEMPR67[31] ), .Y(OR4_70_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%43%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R43C0 (.A_DOUT({
        nc672, nc673, nc674, nc675, nc676,int_R_DATA_TEMPR43[31] , 
       int_R_DATA_TEMPR43[30] ,int_R_DATA_TEMPR43[29] , 
       int_R_DATA_TEMPR43[28] ,int_R_DATA_TEMPR43[27] , 
       int_R_DATA_TEMPR43[26] ,int_R_DATA_TEMPR43[25] , 
       int_R_DATA_TEMPR43[24] ,int_R_DATA_TEMPR43[23] , 
       int_R_DATA_TEMPR43[22] ,int_R_DATA_TEMPR43[21] , 
       int_R_DATA_TEMPR43[20] ,int_R_DATA_TEMPR43[19] , 
       int_R_DATA_TEMPR43[18] ,int_R_DATA_TEMPR43[17] }), .B_DOUT({nc677, 
        nc678, nc679,int_R_DATA_TEMPR43[16] ,int_R_DATA_TEMPR43[15] , 
       int_R_DATA_TEMPR43[14] ,int_R_DATA_TEMPR43[13] , 
       int_R_DATA_TEMPR43[12] ,int_R_DATA_TEMPR43[11] , 
       int_R_DATA_TEMPR43[10] ,int_R_DATA_TEMPR43[9] ,int_R_DATA_TEMPR43[8] , 
       int_R_DATA_TEMPR43[7] ,int_R_DATA_TEMPR43[6] ,int_R_DATA_TEMPR43[5] , 
       int_R_DATA_TEMPR43[4] ,int_R_DATA_TEMPR43[3] ,int_R_DATA_TEMPR43[2] , 
       int_R_DATA_TEMPR43[1] ,int_R_DATA_TEMPR43[0] }), .DB_DETECT( int_DB_DETECT_NG[43] ), .SB_CORRECT(int_SB_CORRECT_NG[43] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[43] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[10] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[10] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_588 (.A(sel_R_DATA_TEMPR40[14] ), .B(sel_R_DATA_TEMPR41[14] ), 
        .C(sel_R_DATA_TEMPR42[14] ), .D(sel_R_DATA_TEMPR43[14] ), .Y(
        OR4_588_Y));
    OR4 OR4_58 (.A(sel_R_DATA_TEMPR40[2] ), .B(sel_R_DATA_TEMPR41[2] ), .C(sel_R_DATA_TEMPR42[2] ), .D(sel_R_DATA_TEMPR43[2] ), .Y(OR4_58_Y));
    OR4 OR4_1112 (.A(sel_R_DATA_TEMPR8[17] ), .B(sel_R_DATA_TEMPR9[17] ), .C(sel_R_DATA_TEMPR10[17] ), .D(sel_R_DATA_TEMPR11[17] ), .Y(OR4_1112_Y)
        );
    AND4 \AND4DB_DETECT[25]  (.A(sel_DB_DETECT_NG[25] ), .B(
        \BLKY2_pipe[6] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[25] ));
    OR4 OR4_276 (.A(sel_R_DATA_TEMPR48[14] ), .B(sel_R_DATA_TEMPR49[14] ), 
        .C(sel_R_DATA_TEMPR50[14] ), .D(sel_R_DATA_TEMPR51[14] ), .Y(
        OR4_276_Y));
    OR4 OR4_242 (.A(sel_R_DATA_TEMPR88[0] ), .B(sel_R_DATA_TEMPR89[0] ), .C(sel_R_DATA_TEMPR90[0] ), .D(sel_R_DATA_TEMPR91[0] ), .Y(OR4_242_Y));
    OR4 OR4_77 (.A(OR4_748_Y), .B(OR4_579_Y), .C(OR4_289_Y), .D(
        OR4_132_Y), .Y(OR4_77_Y));
    OR4 OR4_1370 (.A(sel_R_DATA_TEMPR72[0] ), .B(sel_R_DATA_TEMPR73[0] ), .C(sel_R_DATA_TEMPR74[0] ), .D(sel_R_DATA_TEMPR75[0] ), .Y(OR4_1370_Y));
    OR4 OR4_1354 (.A(sel_R_DATA_TEMPR68[11] ), .B(sel_R_DATA_TEMPR69[11] ), 
        .C(sel_R_DATA_TEMPR70[11] ), .D(sel_R_DATA_TEMPR71[11] ), .Y(
        OR4_1354_Y));
    AND4 \AND4SB_CORRECT[54]  (.A(sel_SB_CORRECT_NG[54] ), .B(
        \BLKY2_pipe[13] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[54] ));
    OR4 OR4_604 (.A(sel_R_DATA_TEMPR52[6] ), .B(sel_R_DATA_TEMPR53[6] ), .C(sel_R_DATA_TEMPR54[6] ), .D(sel_R_DATA_TEMPR55[6] ), .Y(OR4_604_Y));
    OR4 OR4_1124 (.A(sel_R_DATA_TEMPR76[15] ), .B(sel_R_DATA_TEMPR77[15] ), 
        .C(sel_R_DATA_TEMPR78[15] ), .D(sel_R_DATA_TEMPR79[15] ), .Y(
        OR4_1124_Y));
    OR4 OR4_299 (.A(OR4_408_Y), .B(OR4_1177_Y), .C(OR4_321_Y), .D(
        OR4_972_Y), .Y(OR4_299_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[16]  (.A(CFG3_13_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[16] ));
    OR4 OR4_1094 (.A(OR4_29_Y), .B(OR4_749_Y), .C(OR4_47_Y), .D(
        OR4_269_Y), .Y(OR4_1094_Y));
    OR4 OR4_1101 (.A(sel_R_DATA_TEMPR72[3] ), .B(sel_R_DATA_TEMPR73[3] ), .C(sel_R_DATA_TEMPR74[3] ), .D(sel_R_DATA_TEMPR75[3] ), .Y(OR4_1101_Y));
    OR4 OR4_674 (.A(\DB_DETECT[72] ), .B(\DB_DETECT[73] ), .C(
        \DB_DETECT[74] ), .D(\DB_DETECT[75] ), .Y(OR4_674_Y));
    OR4 OR4_455 (.A(sel_R_DATA_TEMPR44[10] ), .B(sel_R_DATA_TEMPR45[10] ), 
        .C(sel_R_DATA_TEMPR46[10] ), .D(sel_R_DATA_TEMPR47[10] ), .Y(
        OR4_455_Y));
    OR4 OR4_486 (.A(OR4_233_Y), .B(OR4_1355_Y), .C(OR4_1326_Y), .D(
        OR4_589_Y), .Y(OR4_486_Y));
    OR4 OR4_1393 (.A(OR4_67_Y), .B(OR4_1288_Y), .C(OR4_964_Y), .D(
        OR4_825_Y), .Y(OR4_1393_Y));
    OR4 \OR4_R_DATA[5]  (.A(OR4_223_Y), .B(OR4_1319_Y), .C(OR4_866_Y), 
        .D(OR4_1146_Y), .Y(R_DATA[5]));
    AND4 \AND4DB_DETECT[52]  (.A(sel_DB_DETECT_NG[52] ), .B(
        \BLKY2_pipe[13] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[52] ));
    OR4 OR4_340 (.A(sel_R_DATA_TEMPR12[29] ), .B(sel_R_DATA_TEMPR13[29] ), 
        .C(sel_R_DATA_TEMPR14[29] ), .D(sel_R_DATA_TEMPR15[29] ), .Y(
        OR4_340_Y));
    OR4 OR4_1066 (.A(sel_R_DATA_TEMPR92[18] ), .B(sel_R_DATA_TEMPR93[18] ), 
        .C(sel_R_DATA_TEMPR94[18] ), .D(sel_R_DATA_TEMPR95[18] ), .Y(
        OR4_1066_Y));
    OR4 OR4_1135 (.A(sel_R_DATA_TEMPR28[18] ), .B(sel_R_DATA_TEMPR29[18] ), 
        .C(sel_R_DATA_TEMPR30[18] ), .D(sel_R_DATA_TEMPR31[18] ), .Y(
        OR4_1135_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[24]  (.D(\BLKY2[24] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[24] ));
    OR4 OR4_719 (.A(sel_R_DATA_TEMPR60[25] ), .B(sel_R_DATA_TEMPR61[25] ), 
        .C(sel_R_DATA_TEMPR62[25] ), .D(sel_R_DATA_TEMPR63[25] ), .Y(
        OR4_719_Y));
    OR4 OR4_1228 (.A(sel_R_DATA_TEMPR68[22] ), .B(sel_R_DATA_TEMPR69[22] ), 
        .C(sel_R_DATA_TEMPR70[22] ), .D(sel_R_DATA_TEMPR71[22] ), .Y(
        OR4_1228_Y));
    OR4 OR4_820 (.A(sel_R_DATA_TEMPR36[9] ), .B(sel_R_DATA_TEMPR37[9] ), .C(sel_R_DATA_TEMPR38[9] ), .D(sel_R_DATA_TEMPR39[9] ), .Y(OR4_820_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%10%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R10C0 (.A_DOUT({
        nc680, nc681, nc682, nc683, nc684,int_R_DATA_TEMPR10[31] , 
       int_R_DATA_TEMPR10[30] ,int_R_DATA_TEMPR10[29] , 
       int_R_DATA_TEMPR10[28] ,int_R_DATA_TEMPR10[27] , 
       int_R_DATA_TEMPR10[26] ,int_R_DATA_TEMPR10[25] , 
       int_R_DATA_TEMPR10[24] ,int_R_DATA_TEMPR10[23] , 
       int_R_DATA_TEMPR10[22] ,int_R_DATA_TEMPR10[21] , 
       int_R_DATA_TEMPR10[20] ,int_R_DATA_TEMPR10[19] , 
       int_R_DATA_TEMPR10[18] ,int_R_DATA_TEMPR10[17] }), .B_DOUT({nc685, 
        nc686, nc687,int_R_DATA_TEMPR10[16] ,int_R_DATA_TEMPR10[15] , 
       int_R_DATA_TEMPR10[14] ,int_R_DATA_TEMPR10[13] , 
       int_R_DATA_TEMPR10[12] ,int_R_DATA_TEMPR10[11] , 
       int_R_DATA_TEMPR10[10] ,int_R_DATA_TEMPR10[9] ,int_R_DATA_TEMPR10[8] , 
       int_R_DATA_TEMPR10[7] ,int_R_DATA_TEMPR10[6] ,int_R_DATA_TEMPR10[5] , 
       int_R_DATA_TEMPR10[4] ,int_R_DATA_TEMPR10[3] ,int_R_DATA_TEMPR10[2] , 
       int_R_DATA_TEMPR10[1] ,int_R_DATA_TEMPR10[0] }), .DB_DETECT( int_DB_DETECT_NG[10] ), .SB_CORRECT(int_SB_CORRECT_NG[10] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[10] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[2] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1031 (.A(OR4_794_Y), .B(OR4_1021_Y), .C(OR4_1193_Y), .D(
        OR4_871_Y), .Y(OR4_1031_Y));
    OR4 OR4_899 (.A(OR4_88_Y), .B(OR4_943_Y), .C(OR4_1163_Y), .D(
        OR4_270_Y), .Y(OR4_899_Y));
    AND4 \AND4SB_CORRECT[102]  (.A(sel_SB_CORRECT_NG[102] ), .B(
        \BLKY2_pipe[25] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[102] ));
    OR4 \OR4_R_DATA[11]  (.A(OR4_2_Y), .B(OR4_1325_Y), .C(OR4_1353_Y), 
        .D(OR4_913_Y), .Y(R_DATA[11]));
    OR4 OR4_122 (.A(sel_R_DATA_TEMPR52[2] ), .B(sel_R_DATA_TEMPR53[2] ), .C(sel_R_DATA_TEMPR54[2] ), .D(sel_R_DATA_TEMPR55[2] ), .Y(OR4_122_Y));
    OR4 OR4_1361 (.A(OR4_12_Y), .B(OR4_432_Y), .C(OR4_102_Y), .D(
        OR4_155_Y), .Y(OR4_1361_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[18]  (.D(\BLKY2[18] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[18] ));
    OR4 OR4_843 (.A(sel_R_DATA_TEMPR104[2] ), .B(sel_R_DATA_TEMPR105[2] ), 
        .C(sel_R_DATA_TEMPR106[2] ), .D(sel_R_DATA_TEMPR107[2] ), .Y(
        OR4_843_Y));
    OR4 OR4_814 (.A(OR4_1025_Y), .B(OR4_1258_Y), .C(OR4_14_Y), .D(
        OR4_755_Y), .Y(OR4_814_Y));
    OR4 OR4_382 (.A(sel_R_DATA_TEMPR116[24] ), .B(sel_R_DATA_TEMPR117[24] ), 
        .C(sel_R_DATA_TEMPR118[24] ), .D(sel_R_DATA_TEMPR119[24] ), .Y(
        OR4_382_Y));
    OR4 OR4_925 (.A(sel_R_DATA_TEMPR32[9] ), .B(sel_R_DATA_TEMPR33[9] ), .C(sel_R_DATA_TEMPR34[9] ), .D(sel_R_DATA_TEMPR35[9] ), .Y(OR4_925_Y));
    OR4 \OR4_R_DATA[9]  (.A(OR4_181_Y), .B(OR4_449_Y), .C(OR4_787_Y), 
        .D(OR4_1061_Y), .Y(R_DATA[9]));
    OR4 OR4_1359 (.A(sel_R_DATA_TEMPR112[15] ), .B(sel_R_DATA_TEMPR113[15] ), 
        .C(sel_R_DATA_TEMPR114[15] ), .D(sel_R_DATA_TEMPR115[15] ), .Y(
        OR4_1359_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%108%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R108C0 (.A_DOUT({
        nc688, nc689, nc690, nc691, nc692,int_R_DATA_TEMPR108[31] , 
       int_R_DATA_TEMPR108[30] ,int_R_DATA_TEMPR108[29] , 
       int_R_DATA_TEMPR108[28] ,int_R_DATA_TEMPR108[27] , 
       int_R_DATA_TEMPR108[26] ,int_R_DATA_TEMPR108[25] , 
       int_R_DATA_TEMPR108[24] ,int_R_DATA_TEMPR108[23] , 
       int_R_DATA_TEMPR108[22] ,int_R_DATA_TEMPR108[21] , 
       int_R_DATA_TEMPR108[20] ,int_R_DATA_TEMPR108[19] , 
       int_R_DATA_TEMPR108[18] ,int_R_DATA_TEMPR108[17] }), .B_DOUT({nc693, 
        nc694, nc695,int_R_DATA_TEMPR108[16] ,int_R_DATA_TEMPR108[15] , 
       int_R_DATA_TEMPR108[14] ,int_R_DATA_TEMPR108[13] , 
       int_R_DATA_TEMPR108[12] ,int_R_DATA_TEMPR108[11] , 
       int_R_DATA_TEMPR108[10] ,int_R_DATA_TEMPR108[9] , 
       int_R_DATA_TEMPR108[8] ,int_R_DATA_TEMPR108[7] , 
       int_R_DATA_TEMPR108[6] ,int_R_DATA_TEMPR108[5] , 
       int_R_DATA_TEMPR108[4] ,int_R_DATA_TEMPR108[3] , 
       int_R_DATA_TEMPR108[2] ,int_R_DATA_TEMPR108[1] , 
       int_R_DATA_TEMPR108[0] }), .DB_DETECT(int_DB_DETECT_NG[108] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[108] ), .ACCESS_BUSY(
        ACCESS_BUSY[108] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[27] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[27] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_18 (.A(sel_R_DATA_TEMPR24[1] ), .B(sel_R_DATA_TEMPR25[1] ), .C(sel_R_DATA_TEMPR26[1] ), .D(sel_R_DATA_TEMPR27[1] ), .Y(OR4_18_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%99%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R99C0 (.A_DOUT({
        nc696, nc697, nc698, nc699, nc700,int_R_DATA_TEMPR99[31] , 
       int_R_DATA_TEMPR99[30] ,int_R_DATA_TEMPR99[29] , 
       int_R_DATA_TEMPR99[28] ,int_R_DATA_TEMPR99[27] , 
       int_R_DATA_TEMPR99[26] ,int_R_DATA_TEMPR99[25] , 
       int_R_DATA_TEMPR99[24] ,int_R_DATA_TEMPR99[23] , 
       int_R_DATA_TEMPR99[22] ,int_R_DATA_TEMPR99[21] , 
       int_R_DATA_TEMPR99[20] ,int_R_DATA_TEMPR99[19] , 
       int_R_DATA_TEMPR99[18] ,int_R_DATA_TEMPR99[17] }), .B_DOUT({nc701, 
        nc702, nc703,int_R_DATA_TEMPR99[16] ,int_R_DATA_TEMPR99[15] , 
       int_R_DATA_TEMPR99[14] ,int_R_DATA_TEMPR99[13] , 
       int_R_DATA_TEMPR99[12] ,int_R_DATA_TEMPR99[11] , 
       int_R_DATA_TEMPR99[10] ,int_R_DATA_TEMPR99[9] ,int_R_DATA_TEMPR99[8] , 
       int_R_DATA_TEMPR99[7] ,int_R_DATA_TEMPR99[6] ,int_R_DATA_TEMPR99[5] , 
       int_R_DATA_TEMPR99[4] ,int_R_DATA_TEMPR99[3] ,int_R_DATA_TEMPR99[2] , 
       int_R_DATA_TEMPR99[1] ,int_R_DATA_TEMPR99[0] }), .DB_DETECT( int_DB_DETECT_NG[99] ), .SB_CORRECT(int_SB_CORRECT_NG[99] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[99] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[24] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[24] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_513 (.A(OR4_984_Y), .B(OR4_1264_Y), .C(OR4_778_Y), .D(
        OR4_116_Y), .Y(OR4_513_Y));
    OR4 OR4_34 (.A(OR4_1037_Y), .B(OR4_1063_Y), .C(OR4_135_Y), .D(
        OR4_1006_Y), .Y(OR4_34_Y));
    OR4 OR4_1181 (.A(sel_R_DATA_TEMPR0[2] ), .B(sel_R_DATA_TEMPR1[2] ), .C(sel_R_DATA_TEMPR2[2] ), .D(sel_R_DATA_TEMPR3[2] ), .Y(OR4_1181_Y));
    OR4 OR4_1050 (.A(sel_R_DATA_TEMPR92[9] ), .B(sel_R_DATA_TEMPR93[9] ), .C(sel_R_DATA_TEMPR94[9] ), .D(sel_R_DATA_TEMPR95[9] ), .Y(OR4_1050_Y));
    OR4 OR4_1147 (.A(\SB_CORRECT[68] ), .B(\SB_CORRECT[69] ), .C(
        \SB_CORRECT[70] ), .D(\SB_CORRECT[71] ), .Y(OR4_1147_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[27]  (.D(\BLKY2[27] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[27] ));
    OR4 OR4_1275 (.A(\SB_CORRECT[16] ), .B(\SB_CORRECT[17] ), .C(
        \SB_CORRECT[18] ), .D(\SB_CORRECT[19] ), .Y(OR4_1275_Y));
    OR4 OR4_868 (.A(sel_R_DATA_TEMPR16[26] ), .B(sel_R_DATA_TEMPR17[26] ), 
        .C(sel_R_DATA_TEMPR18[26] ), .D(sel_R_DATA_TEMPR19[26] ), .Y(
        OR4_868_Y));
    AND4 \AND4DB_DETECT[84]  (.A(sel_DB_DETECT_NG[84] ), .B(
        \BLKY2_pipe[21] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[84] ));
    OR4 OR4_454 (.A(sel_R_DATA_TEMPR112[3] ), .B(sel_R_DATA_TEMPR113[3] ), 
        .C(sel_R_DATA_TEMPR114[3] ), .D(sel_R_DATA_TEMPR115[3] ), .Y(
        OR4_454_Y));
    OR4 OR4_1033 (.A(OR4_172_Y), .B(OR4_1200_Y), .C(OR4_1172_Y), .D(
        OR4_455_Y), .Y(OR4_1033_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[11]  (.A(CFG3_19_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[11] ));
    OR4 OR4_1005 (.A(sel_R_DATA_TEMPR56[1] ), .B(sel_R_DATA_TEMPR57[1] ), .C(sel_R_DATA_TEMPR58[1] ), .D(sel_R_DATA_TEMPR59[1] ), .Y(OR4_1005_Y));
    OR4 \OR4_R_DATA[10]  (.A(OR4_1131_Y), .B(OR4_64_Y), .C(OR4_682_Y), 
        .D(OR4_154_Y), .Y(R_DATA[10]));
    AND4 \AND4SB_CORRECT[97]  (.A(sel_SB_CORRECT_NG[97] ), .B(
        \BLKY2_pipe[24] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[97] ));
    OR4 OR4_229 (.A(sel_R_DATA_TEMPR100[15] ), .B(sel_R_DATA_TEMPR101[15] ), 
        .C(sel_R_DATA_TEMPR102[15] ), .D(sel_R_DATA_TEMPR103[15] ), .Y(
        OR4_229_Y));
    AND4 \AND4SB_CORRECT[12]  (.A(sel_SB_CORRECT_NG[12] ), .B(
        \BLKY2_pipe[3] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[12] ));
    OR4 OR4_356 (.A(OR4_139_Y), .B(OR4_630_Y), .C(OR4_1302_Y), .D(
        OR4_127_Y), .Y(OR4_356_Y));
    AND4 \AND4SB_CORRECT[125]  (.A(sel_SB_CORRECT_NG[125] ), .B(
        \BLKY2_pipe[31] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[125] ));
    OR4 OR4_797 (.A(sel_R_DATA_TEMPR24[29] ), .B(sel_R_DATA_TEMPR25[29] ), 
        .C(sel_R_DATA_TEMPR26[29] ), .D(sel_R_DATA_TEMPR27[29] ), .Y(
        OR4_797_Y));
    AND4 \AND4DB_DETECT[77]  (.A(sel_DB_DETECT_NG[77] ), .B(
        \BLKY2_pipe[19] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[77] ));
    OR4 OR4_794 (.A(sel_R_DATA_TEMPR112[8] ), .B(sel_R_DATA_TEMPR113[8] ), 
        .C(sel_R_DATA_TEMPR114[8] ), .D(sel_R_DATA_TEMPR115[8] ), .Y(
        OR4_794_Y));
    OR4 OR4_1096 (.A(sel_R_DATA_TEMPR16[13] ), .B(sel_R_DATA_TEMPR17[13] ), 
        .C(sel_R_DATA_TEMPR18[13] ), .D(sel_R_DATA_TEMPR19[13] ), .Y(
        OR4_1096_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%33%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R33C0 (.A_DOUT({
        nc704, nc705, nc706, nc707, nc708,int_R_DATA_TEMPR33[31] , 
       int_R_DATA_TEMPR33[30] ,int_R_DATA_TEMPR33[29] , 
       int_R_DATA_TEMPR33[28] ,int_R_DATA_TEMPR33[27] , 
       int_R_DATA_TEMPR33[26] ,int_R_DATA_TEMPR33[25] , 
       int_R_DATA_TEMPR33[24] ,int_R_DATA_TEMPR33[23] , 
       int_R_DATA_TEMPR33[22] ,int_R_DATA_TEMPR33[21] , 
       int_R_DATA_TEMPR33[20] ,int_R_DATA_TEMPR33[19] , 
       int_R_DATA_TEMPR33[18] ,int_R_DATA_TEMPR33[17] }), .B_DOUT({nc709, 
        nc710, nc711,int_R_DATA_TEMPR33[16] ,int_R_DATA_TEMPR33[15] , 
       int_R_DATA_TEMPR33[14] ,int_R_DATA_TEMPR33[13] , 
       int_R_DATA_TEMPR33[12] ,int_R_DATA_TEMPR33[11] , 
       int_R_DATA_TEMPR33[10] ,int_R_DATA_TEMPR33[9] ,int_R_DATA_TEMPR33[8] , 
       int_R_DATA_TEMPR33[7] ,int_R_DATA_TEMPR33[6] ,int_R_DATA_TEMPR33[5] , 
       int_R_DATA_TEMPR33[4] ,int_R_DATA_TEMPR33[3] ,int_R_DATA_TEMPR33[2] , 
       int_R_DATA_TEMPR33[1] ,int_R_DATA_TEMPR33[0] }), .DB_DETECT( int_DB_DETECT_NG[33] ), .SB_CORRECT(int_SB_CORRECT_NG[33] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[33] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[8] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[8] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%72%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R72C0 (.A_DOUT({
        nc712, nc713, nc714, nc715, nc716,int_R_DATA_TEMPR72[31] , 
       int_R_DATA_TEMPR72[30] ,int_R_DATA_TEMPR72[29] , 
       int_R_DATA_TEMPR72[28] ,int_R_DATA_TEMPR72[27] , 
       int_R_DATA_TEMPR72[26] ,int_R_DATA_TEMPR72[25] , 
       int_R_DATA_TEMPR72[24] ,int_R_DATA_TEMPR72[23] , 
       int_R_DATA_TEMPR72[22] ,int_R_DATA_TEMPR72[21] , 
       int_R_DATA_TEMPR72[20] ,int_R_DATA_TEMPR72[19] , 
       int_R_DATA_TEMPR72[18] ,int_R_DATA_TEMPR72[17] }), .B_DOUT({nc717, 
        nc718, nc719,int_R_DATA_TEMPR72[16] ,int_R_DATA_TEMPR72[15] , 
       int_R_DATA_TEMPR72[14] ,int_R_DATA_TEMPR72[13] , 
       int_R_DATA_TEMPR72[12] ,int_R_DATA_TEMPR72[11] , 
       int_R_DATA_TEMPR72[10] ,int_R_DATA_TEMPR72[9] ,int_R_DATA_TEMPR72[8] , 
       int_R_DATA_TEMPR72[7] ,int_R_DATA_TEMPR72[6] ,int_R_DATA_TEMPR72[5] , 
       int_R_DATA_TEMPR72[4] ,int_R_DATA_TEMPR72[3] ,int_R_DATA_TEMPR72[2] , 
       int_R_DATA_TEMPR72[1] ,int_R_DATA_TEMPR72[0] }), .DB_DETECT( int_DB_DETECT_NG[72] ), .SB_CORRECT(int_SB_CORRECT_NG[72] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[72] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[18] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[18] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR2 OR2_23 (.A(sel_R_DATA_TEMPR84[27] ), .B(sel_R_DATA_TEMPR85[27] ), .Y(
        OR2_23_Y));
    OR4 OR4_261 (.A(OR4_653_Y), .B(OR4_670_Y), .C(OR4_654_Y), .D(
        OR4_390_Y), .Y(OR4_261_Y));
    OR4 OR4_29 (.A(sel_R_DATA_TEMPR16[5] ), .B(sel_R_DATA_TEMPR17[5] ), .C(sel_R_DATA_TEMPR18[5] ), .D(sel_R_DATA_TEMPR19[5] ), .Y(OR4_29_Y));
    OR4 \OR4_R_DATA[16]  (.A(OR4_642_Y), .B(OR4_9_Y), .C(OR4_266_Y), 
        .D(OR4_329_Y), .Y(R_DATA[16]));
    OR4 OR4_1125 (.A(sel_R_DATA_TEMPR72[15] ), .B(sel_R_DATA_TEMPR73[15] ), 
        .C(sel_R_DATA_TEMPR74[15] ), .D(sel_R_DATA_TEMPR75[15] ), .Y(
        OR4_1125_Y));
    OR4 OR4_280 (.A(OR4_159_Y), .B(OR4_380_Y), .C(OR4_535_Y), .D(
        OR4_281_Y), .Y(OR4_280_Y));
    OR4 OR4_891 (.A(sel_R_DATA_TEMPR36[0] ), .B(sel_R_DATA_TEMPR37[0] ), .C(sel_R_DATA_TEMPR38[0] ), .D(sel_R_DATA_TEMPR39[0] ), .Y(OR4_891_Y));
    OR4 OR4_587 (.A(sel_R_DATA_TEMPR64[27] ), .B(sel_R_DATA_TEMPR65[27] ), 
        .C(sel_R_DATA_TEMPR66[27] ), .D(sel_R_DATA_TEMPR67[27] ), .Y(
        OR4_587_Y));
    OR4 OR4_1021 (.A(sel_R_DATA_TEMPR116[8] ), .B(sel_R_DATA_TEMPR117[8] ), 
        .C(sel_R_DATA_TEMPR118[8] ), .D(sel_R_DATA_TEMPR119[8] ), .Y(
        OR4_1021_Y));
    AND4 \AND4SB_CORRECT[20]  (.A(sel_SB_CORRECT_NG[20] ), .B(
        \BLKY2_pipe[5] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[20] ));
    OR4 OR4_1391 (.A(OR4_1220_Y), .B(OR2_21_Y), .C(sel_R_DATA_TEMPR86[29] ), .D(sel_R_DATA_TEMPR87[29] ), .Y(OR4_1391_Y)
        );
    OR4 OR4_545 (.A(sel_R_DATA_TEMPR12[19] ), .B(sel_R_DATA_TEMPR13[19] ), 
        .C(sel_R_DATA_TEMPR14[19] ), .D(sel_R_DATA_TEMPR15[19] ), .Y(
        OR4_545_Y));
    OR4 OR4_233 (.A(OR4_565_Y), .B(OR4_438_Y), .C(OR4_537_Y), .D(
        OR4_874_Y), .Y(OR4_233_Y));
    OR4 OR4_1085 (.A(OR4_1081_Y), .B(OR2_1_Y), .C(sel_R_DATA_TEMPR86[4] ), 
        .D(sel_R_DATA_TEMPR87[4] ), .Y(OR4_1085_Y));
    OR4 OR4_829 (.A(OR4_1173_Y), .B(OR2_4_Y), .C(sel_R_DATA_TEMPR86[7] ), 
        .D(sel_R_DATA_TEMPR87[7] ), .Y(OR4_829_Y));
    OR4 OR4_562 (.A(OR4_458_Y), .B(OR4_659_Y), .C(OR4_250_Y), .D(
        OR4_22_Y), .Y(OR4_562_Y));
    OR4 OR4_689 (.A(sel_R_DATA_TEMPR20[7] ), .B(sel_R_DATA_TEMPR21[7] ), .C(sel_R_DATA_TEMPR22[7] ), .D(sel_R_DATA_TEMPR23[7] ), .Y(OR4_689_Y));
    AND4 \AND4SB_CORRECT[31]  (.A(sel_SB_CORRECT_NG[31] ), .B(
        \BLKY2_pipe[7] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[31] ));
    OR4 OR4_643 (.A(OR4_587_Y), .B(OR4_373_Y), .C(OR4_123_Y), .D(
        OR4_987_Y), .Y(OR4_643_Y));
    OR4 OR4_938 (.A(sel_R_DATA_TEMPR68[3] ), .B(sel_R_DATA_TEMPR69[3] ), .C(sel_R_DATA_TEMPR70[3] ), .D(sel_R_DATA_TEMPR71[3] ), .Y(OR4_938_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[5]  (.D(\BLKY2[5] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[5] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[4]  (.A(CFG3_18_Y), .B(CFG3_2_Y)
        , .Y(\BLKY2[4] ));
    OR4 OR4_1240 (.A(sel_R_DATA_TEMPR72[25] ), .B(sel_R_DATA_TEMPR73[25] ), 
        .C(sel_R_DATA_TEMPR74[25] ), .D(sel_R_DATA_TEMPR75[25] ), .Y(
        OR4_1240_Y));
    OR4 OR4_1023 (.A(OR4_16_Y), .B(OR4_469_Y), .C(OR4_43_Y), .D(
        OR4_998_Y), .Y(OR4_1023_Y));
    AND4 \AND4DB_DETECT[82]  (.A(sel_DB_DETECT_NG[82] ), .B(
        \BLKY2_pipe[20] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[82] ));
    AND4 \AND4SB_CORRECT[101]  (.A(sel_SB_CORRECT_NG[101] ), .B(
        \BLKY2_pipe[25] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[101] ));
    OR4 OR4_286 (.A(OR4_908_Y), .B(OR4_1188_Y), .C(OR4_1390_Y), .D(
        OR4_1233_Y), .Y(OR4_286_Y));
    OR4 OR4_78 (.A(sel_R_DATA_TEMPR48[17] ), .B(sel_R_DATA_TEMPR49[17] ), .C(sel_R_DATA_TEMPR50[17] ), .D(sel_R_DATA_TEMPR51[17] ), .Y(OR4_78_Y));
    OR4 OR4_1038 (.A(sel_R_DATA_TEMPR108[5] ), .B(sel_R_DATA_TEMPR109[5] ), 
        .C(sel_R_DATA_TEMPR110[5] ), .D(sel_R_DATA_TEMPR111[5] ), .Y(
        OR4_1038_Y));
    OR4 OR4_1219 (.A(sel_R_DATA_TEMPR32[3] ), .B(sel_R_DATA_TEMPR33[3] ), .C(sel_R_DATA_TEMPR34[3] ), .D(sel_R_DATA_TEMPR35[3] ), .Y(OR4_1219_Y));
    OR4 \OR4_R_DATA[8]  (.A(OR4_686_Y), .B(OR4_845_Y), .C(OR4_513_Y), 
        .D(OR4_1031_Y), .Y(R_DATA[8]));
    OR4 OR4_808 (.A(\DB_DETECT[80] ), .B(\DB_DETECT[81] ), .C(
        \DB_DETECT[82] ), .D(\DB_DETECT[83] ), .Y(OR4_808_Y));
    OR4 OR4_1162 (.A(sel_R_DATA_TEMPR8[8] ), .B(sel_R_DATA_TEMPR9[8] ), .C(sel_R_DATA_TEMPR10[8] ), .D(sel_R_DATA_TEMPR11[8] ), .Y(OR4_1162_Y));
    AND4 \AND4SB_CORRECT[48]  (.A(sel_SB_CORRECT_NG[48] ), .B(
        \BLKY2_pipe[12] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[48] ));
    OR4 OR4_564 (.A(sel_R_DATA_TEMPR68[24] ), .B(sel_R_DATA_TEMPR69[24] ), 
        .C(sel_R_DATA_TEMPR70[24] ), .D(sel_R_DATA_TEMPR71[24] ), .Y(
        OR4_564_Y));
    OR4 OR4_1342 (.A(sel_R_DATA_TEMPR124[0] ), .B(sel_R_DATA_TEMPR125[0] ), 
        .C(sel_R_DATA_TEMPR126[0] ), .D(sel_R_DATA_TEMPR127[0] ), .Y(
        OR4_1342_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%26%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R26C0 (.A_DOUT({
        nc720, nc721, nc722, nc723, nc724,int_R_DATA_TEMPR26[31] , 
       int_R_DATA_TEMPR26[30] ,int_R_DATA_TEMPR26[29] , 
       int_R_DATA_TEMPR26[28] ,int_R_DATA_TEMPR26[27] , 
       int_R_DATA_TEMPR26[26] ,int_R_DATA_TEMPR26[25] , 
       int_R_DATA_TEMPR26[24] ,int_R_DATA_TEMPR26[23] , 
       int_R_DATA_TEMPR26[22] ,int_R_DATA_TEMPR26[21] , 
       int_R_DATA_TEMPR26[20] ,int_R_DATA_TEMPR26[19] , 
       int_R_DATA_TEMPR26[18] ,int_R_DATA_TEMPR26[17] }), .B_DOUT({nc725, 
        nc726, nc727,int_R_DATA_TEMPR26[16] ,int_R_DATA_TEMPR26[15] , 
       int_R_DATA_TEMPR26[14] ,int_R_DATA_TEMPR26[13] , 
       int_R_DATA_TEMPR26[12] ,int_R_DATA_TEMPR26[11] , 
       int_R_DATA_TEMPR26[10] ,int_R_DATA_TEMPR26[9] ,int_R_DATA_TEMPR26[8] , 
       int_R_DATA_TEMPR26[7] ,int_R_DATA_TEMPR26[6] ,int_R_DATA_TEMPR26[5] , 
       int_R_DATA_TEMPR26[4] ,int_R_DATA_TEMPR26[3] ,int_R_DATA_TEMPR26[2] , 
       int_R_DATA_TEMPR26[1] ,int_R_DATA_TEMPR26[0] }), .DB_DETECT( int_DB_DETECT_NG[26] ), .SB_CORRECT(int_SB_CORRECT_NG[26] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[26] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[6] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_154 (.A(OR4_1281_Y), .B(OR4_1133_Y), .C(OR4_1256_Y), .D(
        OR4_560_Y), .Y(OR4_154_Y));
    OR4 OR4_727 (.A(sel_R_DATA_TEMPR24[20] ), .B(sel_R_DATA_TEMPR25[20] ), 
        .C(sel_R_DATA_TEMPR26[20] ), .D(sel_R_DATA_TEMPR27[20] ), .Y(
        OR4_727_Y));
    OR2 OR2_21 (.A(sel_R_DATA_TEMPR84[29] ), .B(sel_R_DATA_TEMPR85[29] ), .Y(
        OR2_21_Y));
    OR4 OR4_684 (.A(OR4_81_Y), .B(OR4_1324_Y), .C(OR4_42_Y), .D(
        OR4_255_Y), .Y(OR4_684_Y));
    OR4 OR4_1242 (.A(sel_R_DATA_TEMPR76[14] ), .B(sel_R_DATA_TEMPR77[14] ), 
        .C(sel_R_DATA_TEMPR78[14] ), .D(sel_R_DATA_TEMPR79[14] ), .Y(
        OR4_1242_Y));
    OR4 OR4_1100 (.A(sel_R_DATA_TEMPR24[6] ), .B(sel_R_DATA_TEMPR25[6] ), .C(sel_R_DATA_TEMPR26[6] ), .D(sel_R_DATA_TEMPR27[6] ), .Y(OR4_1100_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[16]  (.D(\BLKY2[16] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[16] ));
    OR4 OR4_949 (.A(sel_R_DATA_TEMPR0[15] ), .B(sel_R_DATA_TEMPR1[15] ), .C(sel_R_DATA_TEMPR2[15] ), .D(sel_R_DATA_TEMPR3[15] ), .Y(OR4_949_Y));
    OR4 OR4_940 (.A(sel_R_DATA_TEMPR36[1] ), .B(sel_R_DATA_TEMPR37[1] ), .C(sel_R_DATA_TEMPR38[1] ), .D(sel_R_DATA_TEMPR39[1] ), .Y(OR4_940_Y));
    OR4 OR4_962 (.A(OR4_1065_Y), .B(OR4_1274_Y), .C(OR4_1254_Y), .D(
        OR4_520_Y), .Y(OR4_962_Y));
    AND4 \AND4SB_CORRECT[60]  (.A(sel_SB_CORRECT_NG[60] ), .B(
        \BLKY2_pipe[15] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[60] ));
    OR4 OR4_724 (.A(OR4_1247_Y), .B(OR4_72_Y), .C(OR4_227_Y), .D(
        OR4_1330_Y), .Y(OR4_724_Y));
    OR4 OR4_638 (.A(sel_R_DATA_TEMPR64[18] ), .B(sel_R_DATA_TEMPR65[18] ), 
        .C(sel_R_DATA_TEMPR66[18] ), .D(sel_R_DATA_TEMPR67[18] ), .Y(
        OR4_638_Y));
    OR4 OR4_997 (.A(OR4_582_Y), .B(OR4_931_Y), .C(OR4_897_Y), .D(
        OR4_183_Y), .Y(OR4_997_Y));
    OR4 OR4_878 (.A(sel_R_DATA_TEMPR4[18] ), .B(sel_R_DATA_TEMPR5[18] ), .C(sel_R_DATA_TEMPR6[18] ), .D(sel_R_DATA_TEMPR7[18] ), .Y(OR4_878_Y));
    AND4 \AND4SB_CORRECT[107]  (.A(sel_SB_CORRECT_NG[107] ), .B(
        \BLKY2_pipe[26] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[107] ));
    OR4 OR4_22 (.A(sel_R_DATA_TEMPR28[22] ), .B(sel_R_DATA_TEMPR29[22] ), .C(sel_R_DATA_TEMPR30[22] ), .D(sel_R_DATA_TEMPR31[22] ), .Y(OR4_22_Y));
    AND4 \AND4DB_DETECT[13]  (.A(sel_DB_DETECT_NG[13] ), .B(
        \BLKY2_pipe[3] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[13] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[15]  (.A(CFG3_21_Y), .B(
        CFG3_20_Y), .Y(\BLKY2[15] ));
    OR4 OR4_1151 (.A(sel_R_DATA_TEMPR4[16] ), .B(sel_R_DATA_TEMPR5[16] ), .C(sel_R_DATA_TEMPR6[16] ), .D(sel_R_DATA_TEMPR7[16] ), .Y(OR4_1151_Y));
    OR4 OR4_143 (.A(sel_R_DATA_TEMPR80[2] ), .B(sel_R_DATA_TEMPR81[2] ), .C(sel_R_DATA_TEMPR82[2] ), .D(sel_R_DATA_TEMPR83[2] ), .Y(OR4_143_Y));
    OR4 OR4_953 (.A(sel_R_DATA_TEMPR28[17] ), .B(sel_R_DATA_TEMPR29[17] ), 
        .C(sel_R_DATA_TEMPR30[17] ), .D(sel_R_DATA_TEMPR31[17] ), .Y(
        OR4_953_Y));
    OR4 OR4_632 (.A(sel_R_DATA_TEMPR72[23] ), .B(sel_R_DATA_TEMPR73[23] ), 
        .C(sel_R_DATA_TEMPR74[23] ), .D(sel_R_DATA_TEMPR75[23] ), .Y(
        OR4_632_Y));
    OR4 OR4_213 (.A(sel_R_DATA_TEMPR120[21] ), .B(sel_R_DATA_TEMPR121[21] ), 
        .C(sel_R_DATA_TEMPR122[21] ), .D(sel_R_DATA_TEMPR123[21] ), .Y(
        OR4_213_Y));
    OR4 OR4_1074 (.A(sel_R_DATA_TEMPR76[2] ), .B(sel_R_DATA_TEMPR77[2] ), .C(sel_R_DATA_TEMPR78[2] ), .D(sel_R_DATA_TEMPR79[2] ), .Y(OR4_1074_Y));
    OR4 OR4_821 (.A(sel_R_DATA_TEMPR12[4] ), .B(sel_R_DATA_TEMPR13[4] ), .C(sel_R_DATA_TEMPR14[4] ), .D(sel_R_DATA_TEMPR15[4] ), .Y(OR4_821_Y));
    OR4 OR4_201 (.A(sel_R_DATA_TEMPR20[18] ), .B(sel_R_DATA_TEMPR21[18] ), 
        .C(sel_R_DATA_TEMPR22[18] ), .D(sel_R_DATA_TEMPR23[18] ), .Y(
        OR4_201_Y));
    OR4 OR4_361 (.A(sel_R_DATA_TEMPR104[10] ), .B(sel_R_DATA_TEMPR105[10] ), 
        .C(sel_R_DATA_TEMPR106[10] ), .D(sel_R_DATA_TEMPR107[10] ), .Y(
        OR4_361_Y));
    OR4 OR4_1244 (.A(OR4_1108_Y), .B(OR4_211_Y), .C(OR4_860_Y), .D(
        OR4_1092_Y), .Y(OR4_1244_Y));
    OR4 OR4_1373 (.A(sel_R_DATA_TEMPR52[9] ), .B(sel_R_DATA_TEMPR53[9] ), .C(sel_R_DATA_TEMPR54[9] ), .D(sel_R_DATA_TEMPR55[9] ), .Y(OR4_1373_Y));
    OR4 OR4_856 (.A(OR4_801_Y), .B(OR4_148_Y), .C(OR4_817_Y), .D(
        OR4_1040_Y), .Y(OR4_856_Y));
    OR4 OR4_751 (.A(sel_R_DATA_TEMPR92[12] ), .B(sel_R_DATA_TEMPR93[12] ), 
        .C(sel_R_DATA_TEMPR94[12] ), .D(sel_R_DATA_TEMPR95[12] ), .Y(
        OR4_751_Y));
    OR2 OR2_13 (.A(sel_R_DATA_TEMPR84[14] ), .B(sel_R_DATA_TEMPR85[14] ), .Y(
        OR2_13_Y));
    OR4 OR4_6 (.A(sel_R_DATA_TEMPR116[11] ), .B(sel_R_DATA_TEMPR117[11] ), 
        .C(sel_R_DATA_TEMPR118[11] ), .D(sel_R_DATA_TEMPR119[11] ), .Y(
        OR4_6_Y));
    OR4 OR4_918 (.A(sel_R_DATA_TEMPR96[25] ), .B(sel_R_DATA_TEMPR97[25] ), 
        .C(sel_R_DATA_TEMPR98[25] ), .D(sel_R_DATA_TEMPR99[25] ), .Y(
        OR4_918_Y));
    OR4 OR4_1347 (.A(sel_R_DATA_TEMPR0[21] ), .B(sel_R_DATA_TEMPR1[21] ), .C(sel_R_DATA_TEMPR2[21] ), .D(sel_R_DATA_TEMPR3[21] ), .Y(OR4_1347_Y));
    OR4 OR4_271 (.A(sel_R_DATA_TEMPR64[14] ), .B(sel_R_DATA_TEMPR65[14] ), 
        .C(sel_R_DATA_TEMPR66[14] ), .D(sel_R_DATA_TEMPR67[14] ), .Y(
        OR4_271_Y));
    OR4 OR4_1180 (.A(sel_R_DATA_TEMPR52[3] ), .B(sel_R_DATA_TEMPR53[3] ), .C(sel_R_DATA_TEMPR54[3] ), .D(sel_R_DATA_TEMPR55[3] ), .Y(OR4_1180_Y));
    OR4 OR4_460 (.A(sel_R_DATA_TEMPR52[19] ), .B(sel_R_DATA_TEMPR53[19] ), 
        .C(sel_R_DATA_TEMPR54[19] ), .D(sel_R_DATA_TEMPR55[19] ), .Y(
        OR4_460_Y));
    OR4 OR4_1300 (.A(sel_R_DATA_TEMPR108[13] ), .B(sel_R_DATA_TEMPR109[13] ), 
        .C(sel_R_DATA_TEMPR110[13] ), .D(sel_R_DATA_TEMPR111[13] ), .Y(
        OR4_1300_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%64%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R64C0 (.A_DOUT({
        nc728, nc729, nc730, nc731, nc732,int_R_DATA_TEMPR64[31] , 
       int_R_DATA_TEMPR64[30] ,int_R_DATA_TEMPR64[29] , 
       int_R_DATA_TEMPR64[28] ,int_R_DATA_TEMPR64[27] , 
       int_R_DATA_TEMPR64[26] ,int_R_DATA_TEMPR64[25] , 
       int_R_DATA_TEMPR64[24] ,int_R_DATA_TEMPR64[23] , 
       int_R_DATA_TEMPR64[22] ,int_R_DATA_TEMPR64[21] , 
       int_R_DATA_TEMPR64[20] ,int_R_DATA_TEMPR64[19] , 
       int_R_DATA_TEMPR64[18] ,int_R_DATA_TEMPR64[17] }), .B_DOUT({nc733, 
        nc734, nc735,int_R_DATA_TEMPR64[16] ,int_R_DATA_TEMPR64[15] , 
       int_R_DATA_TEMPR64[14] ,int_R_DATA_TEMPR64[13] , 
       int_R_DATA_TEMPR64[12] ,int_R_DATA_TEMPR64[11] , 
       int_R_DATA_TEMPR64[10] ,int_R_DATA_TEMPR64[9] ,int_R_DATA_TEMPR64[8] , 
       int_R_DATA_TEMPR64[7] ,int_R_DATA_TEMPR64[6] ,int_R_DATA_TEMPR64[5] , 
       int_R_DATA_TEMPR64[4] ,int_R_DATA_TEMPR64[3] ,int_R_DATA_TEMPR64[2] , 
       int_R_DATA_TEMPR64[1] ,int_R_DATA_TEMPR64[0] }), .DB_DETECT( int_DB_DETECT_NG[64] ), .SB_CORRECT(int_SB_CORRECT_NG[64] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[64] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[16] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[16] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1028 (.A(sel_R_DATA_TEMPR68[31] ), .B(sel_R_DATA_TEMPR69[31] ), 
        .C(sel_R_DATA_TEMPR70[31] ), .D(sel_R_DATA_TEMPR71[31] ), .Y(
        OR4_1028_Y));
    AND4 \AND4SB_CORRECT[75]  (.A(sel_SB_CORRECT_NG[75] ), .B(
        \BLKY2_pipe[18] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[75] ));
    AND4 \AND4SB_CORRECT[76]  (.A(sel_SB_CORRECT_NG[76] ), .B(
        \BLKY2_pipe[19] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[76] ));
    OR4 OR4_502 (.A(sel_R_DATA_TEMPR120[27] ), .B(sel_R_DATA_TEMPR121[27] ), 
        .C(sel_R_DATA_TEMPR122[27] ), .D(sel_R_DATA_TEMPR123[27] ), .Y(
        OR4_502_Y));
    OR4 OR4_556 (.A(sel_R_DATA_TEMPR52[31] ), .B(sel_R_DATA_TEMPR53[31] ), 
        .C(sel_R_DATA_TEMPR54[31] ), .D(sel_R_DATA_TEMPR55[31] ), .Y(
        OR4_556_Y));
    OR4 OR4_495 (.A(sel_R_DATA_TEMPR112[25] ), .B(sel_R_DATA_TEMPR113[25] ), 
        .C(sel_R_DATA_TEMPR114[25] ), .D(sel_R_DATA_TEMPR115[25] ), .Y(
        OR4_495_Y));
    OR4 OR4_1192 (.A(OR4_1317_Y), .B(OR4_793_Y), .C(OR4_1295_Y), .D(
        OR4_810_Y), .Y(OR4_1192_Y));
    OR4 OR4_835 (.A(sel_R_DATA_TEMPR116[13] ), .B(sel_R_DATA_TEMPR117[13] ), 
        .C(sel_R_DATA_TEMPR118[13] ), .D(sel_R_DATA_TEMPR119[13] ), .Y(
        OR4_835_Y));
    OR4 OR4_572 (.A(sel_R_DATA_TEMPR108[0] ), .B(sel_R_DATA_TEMPR109[0] ), 
        .C(sel_R_DATA_TEMPR110[0] ), .D(sel_R_DATA_TEMPR111[0] ), .Y(
        OR4_572_Y));
    OR4 OR4_618 (.A(OR4_1359_Y), .B(OR4_1221_Y), .C(OR4_1314_Y), .D(
        OR4_973_Y), .Y(OR4_618_Y));
    OR4 OR4_1055 (.A(OR4_160_Y), .B(OR4_418_Y), .C(OR4_168_Y), .D(
        OR4_875_Y), .Y(OR4_1055_Y));
    OR4 OR4_1037 (.A(sel_R_DATA_TEMPR32[24] ), .B(sel_R_DATA_TEMPR33[24] ), 
        .C(sel_R_DATA_TEMPR34[24] ), .D(sel_R_DATA_TEMPR35[24] ), .Y(
        OR4_1037_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%116%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R116C0 (.A_DOUT({
        nc736, nc737, nc738, nc739, nc740,int_R_DATA_TEMPR116[31] , 
       int_R_DATA_TEMPR116[30] ,int_R_DATA_TEMPR116[29] , 
       int_R_DATA_TEMPR116[28] ,int_R_DATA_TEMPR116[27] , 
       int_R_DATA_TEMPR116[26] ,int_R_DATA_TEMPR116[25] , 
       int_R_DATA_TEMPR116[24] ,int_R_DATA_TEMPR116[23] , 
       int_R_DATA_TEMPR116[22] ,int_R_DATA_TEMPR116[21] , 
       int_R_DATA_TEMPR116[20] ,int_R_DATA_TEMPR116[19] , 
       int_R_DATA_TEMPR116[18] ,int_R_DATA_TEMPR116[17] }), .B_DOUT({nc741, 
        nc742, nc743,int_R_DATA_TEMPR116[16] ,int_R_DATA_TEMPR116[15] , 
       int_R_DATA_TEMPR116[14] ,int_R_DATA_TEMPR116[13] , 
       int_R_DATA_TEMPR116[12] ,int_R_DATA_TEMPR116[11] , 
       int_R_DATA_TEMPR116[10] ,int_R_DATA_TEMPR116[9] , 
       int_R_DATA_TEMPR116[8] ,int_R_DATA_TEMPR116[7] , 
       int_R_DATA_TEMPR116[6] ,int_R_DATA_TEMPR116[5] , 
       int_R_DATA_TEMPR116[4] ,int_R_DATA_TEMPR116[3] , 
       int_R_DATA_TEMPR116[2] ,int_R_DATA_TEMPR116[1] , 
       int_R_DATA_TEMPR116[0] }), .DB_DETECT(int_DB_DETECT_NG[116] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[116] ), .ACCESS_BUSY(
        ACCESS_BUSY[116] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[29] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[29] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%97%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R97C0 (.A_DOUT({
        nc744, nc745, nc746, nc747, nc748,int_R_DATA_TEMPR97[31] , 
       int_R_DATA_TEMPR97[30] ,int_R_DATA_TEMPR97[29] , 
       int_R_DATA_TEMPR97[28] ,int_R_DATA_TEMPR97[27] , 
       int_R_DATA_TEMPR97[26] ,int_R_DATA_TEMPR97[25] , 
       int_R_DATA_TEMPR97[24] ,int_R_DATA_TEMPR97[23] , 
       int_R_DATA_TEMPR97[22] ,int_R_DATA_TEMPR97[21] , 
       int_R_DATA_TEMPR97[20] ,int_R_DATA_TEMPR97[19] , 
       int_R_DATA_TEMPR97[18] ,int_R_DATA_TEMPR97[17] }), .B_DOUT({nc749, 
        nc750, nc751,int_R_DATA_TEMPR97[16] ,int_R_DATA_TEMPR97[15] , 
       int_R_DATA_TEMPR97[14] ,int_R_DATA_TEMPR97[13] , 
       int_R_DATA_TEMPR97[12] ,int_R_DATA_TEMPR97[11] , 
       int_R_DATA_TEMPR97[10] ,int_R_DATA_TEMPR97[9] ,int_R_DATA_TEMPR97[8] , 
       int_R_DATA_TEMPR97[7] ,int_R_DATA_TEMPR97[6] ,int_R_DATA_TEMPR97[5] , 
       int_R_DATA_TEMPR97[4] ,int_R_DATA_TEMPR97[3] ,int_R_DATA_TEMPR97[2] , 
       int_R_DATA_TEMPR97[1] ,int_R_DATA_TEMPR97[0] }), .DB_DETECT( int_DB_DETECT_NG[97] ), .SB_CORRECT(int_SB_CORRECT_NG[97] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[97] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[24] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[24] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    CFG3 #( .INIT(8'h10) )  CFG3_8 (.A(W_ADDR[13]), .B(W_ADDR[12]), .C(
        W_ADDR[11]), .Y(CFG3_8_Y));
    OR4 OR4_840 (.A(sel_R_DATA_TEMPR100[19] ), .B(sel_R_DATA_TEMPR101[19] ), 
        .C(sel_R_DATA_TEMPR102[19] ), .D(sel_R_DATA_TEMPR103[19] ), .Y(
        OR4_840_Y));
    OR4 OR4_927 (.A(sel_R_DATA_TEMPR28[25] ), .B(sel_R_DATA_TEMPR29[25] ), 
        .C(sel_R_DATA_TEMPR30[25] ), .D(sel_R_DATA_TEMPR31[25] ), .Y(
        OR4_927_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[0]  (.A(CFG3_16_Y), .B(CFG3_2_Y)
        , .Y(\BLKY2[0] ));
    OR4 \OR4_R_DATA[17]  (.A(OR4_299_Y), .B(OR4_951_Y), .C(OR4_1311_Y), 
        .D(OR4_54_Y), .Y(R_DATA[17]));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%73%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R73C0 (.A_DOUT({
        nc752, nc753, nc754, nc755, nc756,int_R_DATA_TEMPR73[31] , 
       int_R_DATA_TEMPR73[30] ,int_R_DATA_TEMPR73[29] , 
       int_R_DATA_TEMPR73[28] ,int_R_DATA_TEMPR73[27] , 
       int_R_DATA_TEMPR73[26] ,int_R_DATA_TEMPR73[25] , 
       int_R_DATA_TEMPR73[24] ,int_R_DATA_TEMPR73[23] , 
       int_R_DATA_TEMPR73[22] ,int_R_DATA_TEMPR73[21] , 
       int_R_DATA_TEMPR73[20] ,int_R_DATA_TEMPR73[19] , 
       int_R_DATA_TEMPR73[18] ,int_R_DATA_TEMPR73[17] }), .B_DOUT({nc757, 
        nc758, nc759,int_R_DATA_TEMPR73[16] ,int_R_DATA_TEMPR73[15] , 
       int_R_DATA_TEMPR73[14] ,int_R_DATA_TEMPR73[13] , 
       int_R_DATA_TEMPR73[12] ,int_R_DATA_TEMPR73[11] , 
       int_R_DATA_TEMPR73[10] ,int_R_DATA_TEMPR73[9] ,int_R_DATA_TEMPR73[8] , 
       int_R_DATA_TEMPR73[7] ,int_R_DATA_TEMPR73[6] ,int_R_DATA_TEMPR73[5] , 
       int_R_DATA_TEMPR73[4] ,int_R_DATA_TEMPR73[3] ,int_R_DATA_TEMPR73[2] , 
       int_R_DATA_TEMPR73[1] ,int_R_DATA_TEMPR73[0] }), .DB_DETECT( int_DB_DETECT_NG[73] ), .SB_CORRECT(int_SB_CORRECT_NG[73] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[73] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[18] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[18] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_142 (.A(sel_R_DATA_TEMPR16[30] ), .B(sel_R_DATA_TEMPR17[30] ), 
        .C(sel_R_DATA_TEMPR18[30] ), .D(sel_R_DATA_TEMPR19[30] ), .Y(
        OR4_142_Y));
    OR4 OR4_612 (.A(\DB_DETECT[76] ), .B(\DB_DETECT[77] ), .C(
        \DB_DETECT[78] ), .D(\DB_DETECT[79] ), .Y(OR4_612_Y));
    OR4 OR4_504 (.A(sel_R_DATA_TEMPR0[25] ), .B(sel_R_DATA_TEMPR1[25] ), .C(sel_R_DATA_TEMPR2[25] ), .D(sel_R_DATA_TEMPR3[25] ), .Y(OR4_504_Y));
    OR4 OR4_1380 (.A(sel_R_DATA_TEMPR4[23] ), .B(sel_R_DATA_TEMPR5[23] ), .C(sel_R_DATA_TEMPR6[23] ), .D(sel_R_DATA_TEMPR7[23] ), .Y(OR4_1380_Y));
    OR4 OR4_945 (.A(sel_R_DATA_TEMPR16[8] ), .B(sel_R_DATA_TEMPR17[8] ), .C(sel_R_DATA_TEMPR18[8] ), .D(sel_R_DATA_TEMPR19[8] ), .Y(OR4_945_Y));
    OR4 OR4_902 (.A(sel_R_DATA_TEMPR108[25] ), .B(sel_R_DATA_TEMPR109[25] ), 
        .C(sel_R_DATA_TEMPR110[25] ), .D(sel_R_DATA_TEMPR111[25] ), .Y(
        OR4_902_Y));
    OR4 OR4_1076 (.A(sel_R_DATA_TEMPR124[29] ), .B(sel_R_DATA_TEMPR125[29] ), 
        .C(sel_R_DATA_TEMPR126[29] ), .D(sel_R_DATA_TEMPR127[29] ), .Y(
        OR4_1076_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[17]  (.A(CFG3_8_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[17] ));
    OR4 OR4_574 (.A(sel_R_DATA_TEMPR96[19] ), .B(sel_R_DATA_TEMPR97[19] ), 
        .C(sel_R_DATA_TEMPR98[19] ), .D(sel_R_DATA_TEMPR99[19] ), .Y(
        OR4_574_Y));
    OR2 OR2_11 (.A(sel_R_DATA_TEMPR84[21] ), .B(sel_R_DATA_TEMPR85[21] ), .Y(
        OR2_11_Y));
    OR4 OR4_1205 (.A(sel_R_DATA_TEMPR92[3] ), .B(sel_R_DATA_TEMPR93[3] ), .C(sel_R_DATA_TEMPR94[3] ), .D(sel_R_DATA_TEMPR95[3] ), .Y(OR4_1205_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%12%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R12C0 (.A_DOUT({
        nc760, nc761, nc762, nc763, nc764,int_R_DATA_TEMPR12[31] , 
       int_R_DATA_TEMPR12[30] ,int_R_DATA_TEMPR12[29] , 
       int_R_DATA_TEMPR12[28] ,int_R_DATA_TEMPR12[27] , 
       int_R_DATA_TEMPR12[26] ,int_R_DATA_TEMPR12[25] , 
       int_R_DATA_TEMPR12[24] ,int_R_DATA_TEMPR12[23] , 
       int_R_DATA_TEMPR12[22] ,int_R_DATA_TEMPR12[21] , 
       int_R_DATA_TEMPR12[20] ,int_R_DATA_TEMPR12[19] , 
       int_R_DATA_TEMPR12[18] ,int_R_DATA_TEMPR12[17] }), .B_DOUT({nc765, 
        nc766, nc767,int_R_DATA_TEMPR12[16] ,int_R_DATA_TEMPR12[15] , 
       int_R_DATA_TEMPR12[14] ,int_R_DATA_TEMPR12[13] , 
       int_R_DATA_TEMPR12[12] ,int_R_DATA_TEMPR12[11] , 
       int_R_DATA_TEMPR12[10] ,int_R_DATA_TEMPR12[9] ,int_R_DATA_TEMPR12[8] , 
       int_R_DATA_TEMPR12[7] ,int_R_DATA_TEMPR12[6] ,int_R_DATA_TEMPR12[5] , 
       int_R_DATA_TEMPR12[4] ,int_R_DATA_TEMPR12[3] ,int_R_DATA_TEMPR12[2] , 
       int_R_DATA_TEMPR12[1] ,int_R_DATA_TEMPR12[0] }), .DB_DETECT( int_DB_DETECT_NG[12] ), .SB_CORRECT(int_SB_CORRECT_NG[12] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[12] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_494 (.A(sel_R_DATA_TEMPR68[29] ), .B(sel_R_DATA_TEMPR69[29] ), 
        .C(sel_R_DATA_TEMPR70[29] ), .D(sel_R_DATA_TEMPR71[29] ), .Y(
        OR4_494_Y));
    OR4 OR4_1213 (.A(sel_R_DATA_TEMPR68[0] ), .B(sel_R_DATA_TEMPR69[0] ), .C(sel_R_DATA_TEMPR70[0] ), .D(sel_R_DATA_TEMPR71[0] ), .Y(OR4_1213_Y));
    OR4 OR4_972 (.A(OR4_78_Y), .B(OR4_338_Y), .C(OR4_539_Y), .D(
        OR4_377_Y), .Y(OR4_972_Y));
    AND4 \AND4DB_DETECT[50]  (.A(sel_DB_DETECT_NG[50] ), .B(
        \BLKY2_pipe[12] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[50] ));
    OR4 OR4_558 (.A(sel_R_DATA_TEMPR96[23] ), .B(sel_R_DATA_TEMPR97[23] ), 
        .C(sel_R_DATA_TEMPR98[23] ), .D(sel_R_DATA_TEMPR99[23] ), .Y(
        OR4_558_Y));
    OR4 OR4_55 (.A(sel_R_DATA_TEMPR48[30] ), .B(sel_R_DATA_TEMPR49[30] ), .C(sel_R_DATA_TEMPR50[30] ), .D(sel_R_DATA_TEMPR51[30] ), .Y(OR4_55_Y));
    AND4 \AND4DB_DETECT[23]  (.A(sel_DB_DETECT_NG[23] ), .B(
        \BLKY2_pipe[5] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[23] ));
    OR4 OR4_369 (.A(sel_R_DATA_TEMPR72[16] ), .B(sel_R_DATA_TEMPR73[16] ), 
        .C(sel_R_DATA_TEMPR74[16] ), .D(sel_R_DATA_TEMPR75[16] ), .Y(
        OR4_369_Y));
    OR4 OR4_1371 (.A(sel_R_DATA_TEMPR40[21] ), .B(sel_R_DATA_TEMPR41[21] ), 
        .C(sel_R_DATA_TEMPR42[21] ), .D(sel_R_DATA_TEMPR43[21] ), .Y(
        OR4_1371_Y));
    AND4 \AND4DB_DETECT[122]  (.A(sel_DB_DETECT_NG[122] ), .B(
        \BLKY2_pipe[30] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[122] ));
    OR4 OR4_301 (.A(sel_R_DATA_TEMPR92[7] ), .B(sel_R_DATA_TEMPR93[7] ), .C(sel_R_DATA_TEMPR94[7] ), .D(sel_R_DATA_TEMPR95[7] ), .Y(OR4_301_Y));
    AND4 \AND4SB_CORRECT[55]  (.A(sel_SB_CORRECT_NG[55] ), .B(
        \BLKY2_pipe[13] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[55] ));
    AND4 \AND4SB_CORRECT[56]  (.A(sel_SB_CORRECT_NG[56] ), .B(
        \BLKY2_pipe[14] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[56] ));
    AND4 \AND4SB_CORRECT[93]  (.A(sel_SB_CORRECT_NG[93] ), .B(
        \BLKY2_pipe[23] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[93] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%125%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R125C0 (.A_DOUT({
        nc768, nc769, nc770, nc771, nc772,int_R_DATA_TEMPR125[31] , 
       int_R_DATA_TEMPR125[30] ,int_R_DATA_TEMPR125[29] , 
       int_R_DATA_TEMPR125[28] ,int_R_DATA_TEMPR125[27] , 
       int_R_DATA_TEMPR125[26] ,int_R_DATA_TEMPR125[25] , 
       int_R_DATA_TEMPR125[24] ,int_R_DATA_TEMPR125[23] , 
       int_R_DATA_TEMPR125[22] ,int_R_DATA_TEMPR125[21] , 
       int_R_DATA_TEMPR125[20] ,int_R_DATA_TEMPR125[19] , 
       int_R_DATA_TEMPR125[18] ,int_R_DATA_TEMPR125[17] }), .B_DOUT({nc773, 
        nc774, nc775,int_R_DATA_TEMPR125[16] ,int_R_DATA_TEMPR125[15] , 
       int_R_DATA_TEMPR125[14] ,int_R_DATA_TEMPR125[13] , 
       int_R_DATA_TEMPR125[12] ,int_R_DATA_TEMPR125[11] , 
       int_R_DATA_TEMPR125[10] ,int_R_DATA_TEMPR125[9] , 
       int_R_DATA_TEMPR125[8] ,int_R_DATA_TEMPR125[7] , 
       int_R_DATA_TEMPR125[6] ,int_R_DATA_TEMPR125[5] , 
       int_R_DATA_TEMPR125[4] ,int_R_DATA_TEMPR125[3] , 
       int_R_DATA_TEMPR125[2] ,int_R_DATA_TEMPR125[1] , 
       int_R_DATA_TEMPR125[0] }), .DB_DETECT(int_DB_DETECT_NG[125] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[125] ), .ACCESS_BUSY(
        ACCESS_BUSY[125] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[31] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[31] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_396 (.A(sel_R_DATA_TEMPR0[1] ), .B(sel_R_DATA_TEMPR1[1] ), .C(sel_R_DATA_TEMPR2[1] ), .D(sel_R_DATA_TEMPR3[1] ), .Y(OR4_396_Y));
    AND4 \AND4SB_CORRECT[104]  (.A(sel_SB_CORRECT_NG[104] ), .B(
        \BLKY2_pipe[26] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[104] ));
    OR4 OR4_249 (.A(sel_R_DATA_TEMPR72[29] ), .B(sel_R_DATA_TEMPR73[29] ), 
        .C(sel_R_DATA_TEMPR74[29] ), .D(sel_R_DATA_TEMPR75[29] ), .Y(
        OR4_249_Y));
    AND4 \AND4DB_DETECT[0]  (.A(sel_DB_DETECT_NG[0] ), .B(
        \BLKY2_pipe[0] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[0] ));
    OR4 OR4_425 (.A(sel_R_DATA_TEMPR72[30] ), .B(sel_R_DATA_TEMPR73[30] ), 
        .C(sel_R_DATA_TEMPR74[30] ), .D(sel_R_DATA_TEMPR75[30] ), .Y(
        OR4_425_Y));
    OR4 OR4_371 (.A(sel_R_DATA_TEMPR32[7] ), .B(sel_R_DATA_TEMPR33[7] ), .C(sel_R_DATA_TEMPR34[7] ), .D(sel_R_DATA_TEMPR35[7] ), .Y(OR4_371_Y));
    OR4 OR4_815 (.A(sel_R_DATA_TEMPR4[21] ), .B(sel_R_DATA_TEMPR5[21] ), .C(sel_R_DATA_TEMPR6[21] ), .D(sel_R_DATA_TEMPR7[21] ), .Y(OR4_815_Y));
    OR4 OR4_400 (.A(sel_R_DATA_TEMPR32[1] ), .B(sel_R_DATA_TEMPR33[1] ), .C(sel_R_DATA_TEMPR34[1] ), .D(sel_R_DATA_TEMPR35[1] ), .Y(OR4_400_Y));
    OR4 OR4_636 (.A(OR4_1077_Y), .B(OR4_430_Y), .C(OR4_1100_Y), .D(
        OR4_1322_Y), .Y(OR4_636_Y));
    OR4 OR4_456 (.A(sel_R_DATA_TEMPR16[27] ), .B(sel_R_DATA_TEMPR17[27] ), 
        .C(sel_R_DATA_TEMPR18[27] ), .D(sel_R_DATA_TEMPR19[27] ), .Y(
        OR4_456_Y));
    AND4 \AND4DB_DETECT[94]  (.A(sel_DB_DETECT_NG[94] ), .B(
        \BLKY2_pipe[23] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[94] ));
    OR4 OR4_1027 (.A(sel_R_DATA_TEMPR4[29] ), .B(sel_R_DATA_TEMPR5[29] ), .C(sel_R_DATA_TEMPR6[29] ), .D(sel_R_DATA_TEMPR7[29] ), .Y(OR4_1027_Y));
    OR4 OR4_1346 (.A(sel_R_DATA_TEMPR12[28] ), .B(sel_R_DATA_TEMPR13[28] ), 
        .C(sel_R_DATA_TEMPR14[28] ), .D(sel_R_DATA_TEMPR15[28] ), .Y(
        OR4_1346_Y));
    OR4 OR4_1285 (.A(sel_R_DATA_TEMPR8[18] ), .B(sel_R_DATA_TEMPR9[18] ), .C(sel_R_DATA_TEMPR10[18] ), .D(sel_R_DATA_TEMPR11[18] ), .Y(OR4_1285_Y)
        );
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[5]  (.A(CFG3_11_Y), .B(CFG3_2_Y)
        , .Y(\BLKY2[5] ));
    OR4 OR4_1119 (.A(sel_R_DATA_TEMPR56[18] ), .B(sel_R_DATA_TEMPR57[18] ), 
        .C(sel_R_DATA_TEMPR58[18] ), .D(sel_R_DATA_TEMPR59[18] ), .Y(
        OR4_1119_Y));
    OR4 OR4_1269 (.A(sel_R_DATA_TEMPR104[16] ), .B(sel_R_DATA_TEMPR105[16] ), 
        .C(sel_R_DATA_TEMPR106[16] ), .D(sel_R_DATA_TEMPR107[16] ), .Y(
        OR4_1269_Y));
    OR4 OR4_888 (.A(OR4_226_Y), .B(OR4_878_Y), .C(OR4_1285_Y), .D(
        OR4_158_Y), .Y(OR4_888_Y));
    OR4 OR4_470 (.A(sel_R_DATA_TEMPR4[27] ), .B(sel_R_DATA_TEMPR5[27] ), .C(sel_R_DATA_TEMPR6[27] ), .D(sel_R_DATA_TEMPR7[27] ), .Y(OR4_470_Y));
    AND4 \AND4DB_DETECT[47]  (.A(sel_DB_DETECT_NG[47] ), .B(
        \BLKY2_pipe[11] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[47] ));
    OR4 OR4_849 (.A(sel_R_DATA_TEMPR80[13] ), .B(sel_R_DATA_TEMPR81[13] ), 
        .C(sel_R_DATA_TEMPR82[13] ), .D(sel_R_DATA_TEMPR83[13] ), .Y(
        OR4_849_Y));
    AND4 \AND4DB_DETECT[64]  (.A(sel_DB_DETECT_NG[64] ), .B(
        \BLKY2_pipe[16] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[64] ));
    OR4 OR4_1150 (.A(sel_R_DATA_TEMPR96[12] ), .B(sel_R_DATA_TEMPR97[12] ), 
        .C(sel_R_DATA_TEMPR98[12] ), .D(sel_R_DATA_TEMPR99[12] ), .Y(
        OR4_1150_Y));
    AND4 \AND4SB_CORRECT[94]  (.A(sel_SB_CORRECT_NG[94] ), .B(
        \BLKY2_pipe[23] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[94] ));
    OR4 OR4_352 (.A(sel_R_DATA_TEMPR48[6] ), .B(sel_R_DATA_TEMPR49[6] ), .C(sel_R_DATA_TEMPR50[6] ), .D(sel_R_DATA_TEMPR51[6] ), .Y(OR4_352_Y));
    OR4 OR4_15 (.A(OR4_613_Y), .B(OR4_1391_Y), .C(OR4_462_Y), .D(
        OR4_1333_Y), .Y(OR4_15_Y));
    OR4 OR4_424 (.A(sel_R_DATA_TEMPR112[20] ), .B(sel_R_DATA_TEMPR113[20] ), 
        .C(sel_R_DATA_TEMPR114[20] ), .D(sel_R_DATA_TEMPR115[20] ), .Y(
        OR4_424_Y));
    OR4 OR4_281 (.A(sel_R_DATA_TEMPR76[6] ), .B(sel_R_DATA_TEMPR77[6] ), .C(sel_R_DATA_TEMPR78[6] ), .D(sel_R_DATA_TEMPR79[6] ), .Y(OR4_281_Y));
    AND4 \AND4DB_DETECT[120]  (.A(sel_DB_DETECT_NG[120] ), .B(
        \BLKY2_pipe[30] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[120] ));
    AND4 \AND4DB_DETECT[36]  (.A(sel_DB_DETECT_NG[36] ), .B(
        \BLKY2_pipe[9] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[36] ));
    OR4 OR4_769 (.A(OR4_1156_Y), .B(OR4_635_Y), .C(OR4_837_Y), .D(
        OR4_1346_Y), .Y(OR4_769_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%60%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R60C0 (.A_DOUT({
        nc776, nc777, nc778, nc779, nc780,int_R_DATA_TEMPR60[31] , 
       int_R_DATA_TEMPR60[30] ,int_R_DATA_TEMPR60[29] , 
       int_R_DATA_TEMPR60[28] ,int_R_DATA_TEMPR60[27] , 
       int_R_DATA_TEMPR60[26] ,int_R_DATA_TEMPR60[25] , 
       int_R_DATA_TEMPR60[24] ,int_R_DATA_TEMPR60[23] , 
       int_R_DATA_TEMPR60[22] ,int_R_DATA_TEMPR60[21] , 
       int_R_DATA_TEMPR60[20] ,int_R_DATA_TEMPR60[19] , 
       int_R_DATA_TEMPR60[18] ,int_R_DATA_TEMPR60[17] }), .B_DOUT({nc781, 
        nc782, nc783,int_R_DATA_TEMPR60[16] ,int_R_DATA_TEMPR60[15] , 
       int_R_DATA_TEMPR60[14] ,int_R_DATA_TEMPR60[13] , 
       int_R_DATA_TEMPR60[12] ,int_R_DATA_TEMPR60[11] , 
       int_R_DATA_TEMPR60[10] ,int_R_DATA_TEMPR60[9] ,int_R_DATA_TEMPR60[8] , 
       int_R_DATA_TEMPR60[7] ,int_R_DATA_TEMPR60[6] ,int_R_DATA_TEMPR60[5] , 
       int_R_DATA_TEMPR60[4] ,int_R_DATA_TEMPR60[3] ,int_R_DATA_TEMPR60[2] , 
       int_R_DATA_TEMPR60[1] ,int_R_DATA_TEMPR60[0] }), .DB_DETECT( int_DB_DETECT_NG[60] ), .SB_CORRECT(int_SB_CORRECT_NG[60] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[60] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[15] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[15] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4DB_DETECT[31]  (.A(sel_DB_DETECT_NG[31] ), .B(
        \BLKY2_pipe[7] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[31] ));
    OR4 OR4_1116 (.A(OR4_680_Y), .B(OR4_571_Y), .C(OR4_1035_Y), .D(
        OR4_522_Y), .Y(OR4_1116_Y));
    OR4 OR4_864 (.A(sel_R_DATA_TEMPR124[21] ), .B(sel_R_DATA_TEMPR125[21] ), 
        .C(sel_R_DATA_TEMPR126[21] ), .D(sel_R_DATA_TEMPR127[21] ), .Y(
        OR4_864_Y));
    OR4 OR4_194 (.A(sel_R_DATA_TEMPR8[25] ), .B(sel_R_DATA_TEMPR9[25] ), .C(sel_R_DATA_TEMPR10[25] ), .D(sel_R_DATA_TEMPR11[25] ), .Y(OR4_194_Y));
    OR4 OR4_326 (.A(sel_R_DATA_TEMPR52[24] ), .B(sel_R_DATA_TEMPR53[24] ), 
        .C(sel_R_DATA_TEMPR54[24] ), .D(sel_R_DATA_TEMPR55[24] ), .Y(
        OR4_326_Y));
    AND4 \AND4SB_CORRECT[11]  (.A(sel_SB_CORRECT_NG[11] ), .B(
        \BLKY2_pipe[2] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[11] ));
    OR4 OR4_1237 (.A(sel_R_DATA_TEMPR52[25] ), .B(sel_R_DATA_TEMPR53[25] ), 
        .C(sel_R_DATA_TEMPR54[25] ), .D(sel_R_DATA_TEMPR55[25] ), .Y(
        OR4_1237_Y));
    AND4 \AND4DB_DETECT[7]  (.A(sel_DB_DETECT_NG[7] ), .B(
        \BLKY2_pipe[1] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[7] ));
    AND4 \AND4SB_CORRECT[2]  (.A(sel_SB_CORRECT_NG[2] ), .B(
        \BLKY2_pipe[0] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[2] ));
    OR4 OR4_747 (.A(sel_R_DATA_TEMPR96[31] ), .B(sel_R_DATA_TEMPR97[31] ), 
        .C(sel_R_DATA_TEMPR98[31] ), .D(sel_R_DATA_TEMPR99[31] ), .Y(
        OR4_747_Y));
    OR4 OR4_563 (.A(sel_R_DATA_TEMPR8[4] ), .B(sel_R_DATA_TEMPR9[4] ), .C(sel_R_DATA_TEMPR10[4] ), .D(sel_R_DATA_TEMPR11[4] ), .Y(OR4_563_Y));
    OR4 OR4_93 (.A(sel_R_DATA_TEMPR0[6] ), .B(sel_R_DATA_TEMPR1[6] ), .C(sel_R_DATA_TEMPR2[6] ), .D(sel_R_DATA_TEMPR3[6] ), .Y(OR4_93_Y));
    OR4 OR4_1211 (.A(OR4_966_Y), .B(OR4_1277_Y), .C(OR4_34_Y), .D(
        OR4_1042_Y), .Y(OR4_1211_Y));
    OR4 OR4_744 (.A(sel_R_DATA_TEMPR76[29] ), .B(sel_R_DATA_TEMPR77[29] ), 
        .C(sel_R_DATA_TEMPR78[29] ), .D(sel_R_DATA_TEMPR79[29] ), .Y(
        OR4_744_Y));
    OR4 OR4_1350 (.A(OR4_715_Y), .B(OR4_457_Y), .C(OR4_799_Y), .D(
        OR4_652_Y), .Y(OR4_1350_Y));
    OR4 OR4_616 (.A(sel_R_DATA_TEMPR24[13] ), .B(sel_R_DATA_TEMPR25[13] ), 
        .C(sel_R_DATA_TEMPR26[13] ), .D(sel_R_DATA_TEMPR27[13] ), .Y(
        OR4_616_Y));
    OR4 OR4_309 (.A(sel_R_DATA_TEMPR76[19] ), .B(sel_R_DATA_TEMPR77[19] ), 
        .C(sel_R_DATA_TEMPR78[19] ), .D(sel_R_DATA_TEMPR79[19] ), .Y(
        OR4_309_Y));
    OR4 OR4_1118 (.A(sel_R_DATA_TEMPR96[7] ), .B(sel_R_DATA_TEMPR97[7] ), .C(sel_R_DATA_TEMPR98[7] ), .D(sel_R_DATA_TEMPR99[7] ), .Y(OR4_1118_Y));
    OR4 OR4_582 (.A(sel_R_DATA_TEMPR32[13] ), .B(sel_R_DATA_TEMPR33[13] ), 
        .C(sel_R_DATA_TEMPR34[13] ), .D(sel_R_DATA_TEMPR35[13] ), .Y(
        OR4_582_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%102%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R102C0 (.A_DOUT({
        nc784, nc785, nc786, nc787, nc788,int_R_DATA_TEMPR102[31] , 
       int_R_DATA_TEMPR102[30] ,int_R_DATA_TEMPR102[29] , 
       int_R_DATA_TEMPR102[28] ,int_R_DATA_TEMPR102[27] , 
       int_R_DATA_TEMPR102[26] ,int_R_DATA_TEMPR102[25] , 
       int_R_DATA_TEMPR102[24] ,int_R_DATA_TEMPR102[23] , 
       int_R_DATA_TEMPR102[22] ,int_R_DATA_TEMPR102[21] , 
       int_R_DATA_TEMPR102[20] ,int_R_DATA_TEMPR102[19] , 
       int_R_DATA_TEMPR102[18] ,int_R_DATA_TEMPR102[17] }), .B_DOUT({nc789, 
        nc790, nc791,int_R_DATA_TEMPR102[16] ,int_R_DATA_TEMPR102[15] , 
       int_R_DATA_TEMPR102[14] ,int_R_DATA_TEMPR102[13] , 
       int_R_DATA_TEMPR102[12] ,int_R_DATA_TEMPR102[11] , 
       int_R_DATA_TEMPR102[10] ,int_R_DATA_TEMPR102[9] , 
       int_R_DATA_TEMPR102[8] ,int_R_DATA_TEMPR102[7] , 
       int_R_DATA_TEMPR102[6] ,int_R_DATA_TEMPR102[5] , 
       int_R_DATA_TEMPR102[4] ,int_R_DATA_TEMPR102[3] , 
       int_R_DATA_TEMPR102[2] ,int_R_DATA_TEMPR102[1] , 
       int_R_DATA_TEMPR102[0] }), .DB_DETECT(int_DB_DETECT_NG[102] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[102] ), .ACCESS_BUSY(
        ACCESS_BUSY[102] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[25] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[25] , W_ADDR[10], \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_24 (.A(sel_R_DATA_TEMPR120[25] ), .B(sel_R_DATA_TEMPR121[25] ), 
        .C(sel_R_DATA_TEMPR122[25] ), .D(sel_R_DATA_TEMPR123[25] ), .Y(
        OR4_24_Y));
    OR4 OR4_1299 (.A(OR4_814_Y), .B(OR4_1153_Y), .C(OR4_222_Y), .D(
        OR4_595_Y), .Y(OR4_1299_Y));
    AND4 \AND4SB_CORRECT[112]  (.A(sel_SB_CORRECT_NG[112] ), .B(
        \BLKY2_pipe[28] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[112] ));
    AND4 \AND4SB_CORRECT[47]  (.A(sel_SB_CORRECT_NG[47] ), .B(
        \BLKY2_pipe[11] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[47] ));
    OR4 OR4_993 (.A(sel_R_DATA_TEMPR116[12] ), .B(sel_R_DATA_TEMPR117[12] ), 
        .C(sel_R_DATA_TEMPR118[12] ), .D(sel_R_DATA_TEMPR119[12] ), .Y(
        OR4_993_Y));
    AND4 \AND4DB_DETECT[92]  (.A(sel_DB_DETECT_NG[92] ), .B(
        \BLKY2_pipe[23] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[92] ));
    OR4 OR4_8 (.A(sel_R_DATA_TEMPR44[16] ), .B(sel_R_DATA_TEMPR45[16] ), .C(sel_R_DATA_TEMPR46[16] ), .D(sel_R_DATA_TEMPR47[16] ), .Y(OR4_8_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[7]  (.A(CFG3_21_Y), .B(CFG3_2_Y)
        , .Y(\BLKY2[7] ));
    OR4 OR4_379 (.A(OR4_1267_Y), .B(OR4_122_Y), .C(OR4_1048_Y), .D(
        OR4_391_Y), .Y(OR4_379_Y));
    OR4 OR4_1334 (.A(sel_R_DATA_TEMPR40[27] ), .B(sel_R_DATA_TEMPR41[27] ), 
        .C(sel_R_DATA_TEMPR42[27] ), .D(sel_R_DATA_TEMPR43[27] ), .Y(
        OR4_1334_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%54%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R54C0 (.A_DOUT({
        nc792, nc793, nc794, nc795, nc796,int_R_DATA_TEMPR54[31] , 
       int_R_DATA_TEMPR54[30] ,int_R_DATA_TEMPR54[29] , 
       int_R_DATA_TEMPR54[28] ,int_R_DATA_TEMPR54[27] , 
       int_R_DATA_TEMPR54[26] ,int_R_DATA_TEMPR54[25] , 
       int_R_DATA_TEMPR54[24] ,int_R_DATA_TEMPR54[23] , 
       int_R_DATA_TEMPR54[22] ,int_R_DATA_TEMPR54[21] , 
       int_R_DATA_TEMPR54[20] ,int_R_DATA_TEMPR54[19] , 
       int_R_DATA_TEMPR54[18] ,int_R_DATA_TEMPR54[17] }), .B_DOUT({nc797, 
        nc798, nc799,int_R_DATA_TEMPR54[16] ,int_R_DATA_TEMPR54[15] , 
       int_R_DATA_TEMPR54[14] ,int_R_DATA_TEMPR54[13] , 
       int_R_DATA_TEMPR54[12] ,int_R_DATA_TEMPR54[11] , 
       int_R_DATA_TEMPR54[10] ,int_R_DATA_TEMPR54[9] ,int_R_DATA_TEMPR54[8] , 
       int_R_DATA_TEMPR54[7] ,int_R_DATA_TEMPR54[6] ,int_R_DATA_TEMPR54[5] , 
       int_R_DATA_TEMPR54[4] ,int_R_DATA_TEMPR54[3] ,int_R_DATA_TEMPR54[2] , 
       int_R_DATA_TEMPR54[1] ,int_R_DATA_TEMPR54[0] }), .DB_DETECT( int_DB_DETECT_NG[54] ), .SB_CORRECT(int_SB_CORRECT_NG[54] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[54] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[13] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[13] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1004 (.A(sel_R_DATA_TEMPR16[29] ), .B(sel_R_DATA_TEMPR17[29] ), 
        .C(sel_R_DATA_TEMPR18[29] ), .D(sel_R_DATA_TEMPR19[29] ), .Y(
        OR4_1004_Y));
    OR4 OR4_841 (.A(sel_R_DATA_TEMPR0[24] ), .B(sel_R_DATA_TEMPR1[24] ), .C(sel_R_DATA_TEMPR2[24] ), .D(sel_R_DATA_TEMPR3[24] ), .Y(OR4_841_Y));
    OR4 OR4_250 (.A(sel_R_DATA_TEMPR24[22] ), .B(sel_R_DATA_TEMPR25[22] ), 
        .C(sel_R_DATA_TEMPR26[22] ), .D(sel_R_DATA_TEMPR27[22] ), .Y(
        OR4_250_Y));
    AND4 \AND4DB_DETECT[80]  (.A(sel_DB_DETECT_NG[80] ), .B(
        \BLKY2_pipe[20] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[80] ));
    OR4 OR4_1172 (.A(sel_R_DATA_TEMPR40[10] ), .B(sel_R_DATA_TEMPR41[10] ), 
        .C(sel_R_DATA_TEMPR42[10] ), .D(sel_R_DATA_TEMPR43[10] ), .Y(
        OR4_1172_Y));
    OR4 OR4_557 (.A(sel_R_DATA_TEMPR108[1] ), .B(sel_R_DATA_TEMPR109[1] ), 
        .C(sel_R_DATA_TEMPR110[1] ), .D(sel_R_DATA_TEMPR111[1] ), .Y(
        OR4_557_Y));
    AND4 \AND4DB_DETECT[106]  (.A(sel_DB_DETECT_NG[106] ), .B(
        \BLKY2_pipe[26] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[106] ));
    OR4 OR4_896 (.A(sel_R_DATA_TEMPR104[7] ), .B(sel_R_DATA_TEMPR105[7] ), 
        .C(sel_R_DATA_TEMPR106[7] ), .D(sel_R_DATA_TEMPR107[7] ), .Y(
        OR4_896_Y));
    OR2 OR2_4 (.A(sel_R_DATA_TEMPR84[7] ), .B(sel_R_DATA_TEMPR85[7] ), .Y(
        OR2_4_Y));
    OR4 OR4_334 (.A(sel_R_DATA_TEMPR104[23] ), .B(sel_R_DATA_TEMPR105[23] ), 
        .C(sel_R_DATA_TEMPR106[23] ), .D(sel_R_DATA_TEMPR107[23] ), .Y(
        OR4_334_Y));
    OR4 OR4_791 (.A(sel_R_DATA_TEMPR104[28] ), .B(sel_R_DATA_TEMPR105[28] ), 
        .C(sel_R_DATA_TEMPR106[28] ), .D(sel_R_DATA_TEMPR107[28] ), .Y(
        OR4_791_Y));
    OR4 OR4_1303 (.A(OR4_950_Y), .B(OR4_235_Y), .C(OR4_624_Y), .D(
        OR4_884_Y), .Y(OR4_1303_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%100%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R100C0 (.A_DOUT({
        nc800, nc801, nc802, nc803, nc804,int_R_DATA_TEMPR100[31] , 
       int_R_DATA_TEMPR100[30] ,int_R_DATA_TEMPR100[29] , 
       int_R_DATA_TEMPR100[28] ,int_R_DATA_TEMPR100[27] , 
       int_R_DATA_TEMPR100[26] ,int_R_DATA_TEMPR100[25] , 
       int_R_DATA_TEMPR100[24] ,int_R_DATA_TEMPR100[23] , 
       int_R_DATA_TEMPR100[22] ,int_R_DATA_TEMPR100[21] , 
       int_R_DATA_TEMPR100[20] ,int_R_DATA_TEMPR100[19] , 
       int_R_DATA_TEMPR100[18] ,int_R_DATA_TEMPR100[17] }), .B_DOUT({nc805, 
        nc806, nc807,int_R_DATA_TEMPR100[16] ,int_R_DATA_TEMPR100[15] , 
       int_R_DATA_TEMPR100[14] ,int_R_DATA_TEMPR100[13] , 
       int_R_DATA_TEMPR100[12] ,int_R_DATA_TEMPR100[11] , 
       int_R_DATA_TEMPR100[10] ,int_R_DATA_TEMPR100[9] , 
       int_R_DATA_TEMPR100[8] ,int_R_DATA_TEMPR100[7] , 
       int_R_DATA_TEMPR100[6] ,int_R_DATA_TEMPR100[5] , 
       int_R_DATA_TEMPR100[4] ,int_R_DATA_TEMPR100[3] , 
       int_R_DATA_TEMPR100[2] ,int_R_DATA_TEMPR100[1] , 
       int_R_DATA_TEMPR100[0] }), .DB_DETECT(int_DB_DETECT_NG[100] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[100] ), .ACCESS_BUSY(
        ACCESS_BUSY[100] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[25] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[25] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%103%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R103C0 (.A_DOUT({
        nc808, nc809, nc810, nc811, nc812,int_R_DATA_TEMPR103[31] , 
       int_R_DATA_TEMPR103[30] ,int_R_DATA_TEMPR103[29] , 
       int_R_DATA_TEMPR103[28] ,int_R_DATA_TEMPR103[27] , 
       int_R_DATA_TEMPR103[26] ,int_R_DATA_TEMPR103[25] , 
       int_R_DATA_TEMPR103[24] ,int_R_DATA_TEMPR103[23] , 
       int_R_DATA_TEMPR103[22] ,int_R_DATA_TEMPR103[21] , 
       int_R_DATA_TEMPR103[20] ,int_R_DATA_TEMPR103[19] , 
       int_R_DATA_TEMPR103[18] ,int_R_DATA_TEMPR103[17] }), .B_DOUT({nc813, 
        nc814, nc815,int_R_DATA_TEMPR103[16] ,int_R_DATA_TEMPR103[15] , 
       int_R_DATA_TEMPR103[14] ,int_R_DATA_TEMPR103[13] , 
       int_R_DATA_TEMPR103[12] ,int_R_DATA_TEMPR103[11] , 
       int_R_DATA_TEMPR103[10] ,int_R_DATA_TEMPR103[9] , 
       int_R_DATA_TEMPR103[8] ,int_R_DATA_TEMPR103[7] , 
       int_R_DATA_TEMPR103[6] ,int_R_DATA_TEMPR103[5] , 
       int_R_DATA_TEMPR103[4] ,int_R_DATA_TEMPR103[3] , 
       int_R_DATA_TEMPR103[2] ,int_R_DATA_TEMPR103[1] , 
       int_R_DATA_TEMPR103[0] }), .DB_DETECT(int_DB_DETECT_NG[103] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[103] ), .ACCESS_BUSY(
        ACCESS_BUSY[103] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[25] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[25] , W_ADDR[10], W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4DB_DETECT[62]  (.A(sel_DB_DETECT_NG[62] ), .B(
        \BLKY2_pipe[15] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[62] ));
    OR4 OR4_1144 (.A(sel_R_DATA_TEMPR92[11] ), .B(sel_R_DATA_TEMPR93[11] ), 
        .C(sel_R_DATA_TEMPR94[11] ), .D(sel_R_DATA_TEMPR95[11] ), .Y(
        OR4_1144_Y));
    OR4 OR4_131 (.A(sel_R_DATA_TEMPR12[21] ), .B(sel_R_DATA_TEMPR13[21] ), 
        .C(sel_R_DATA_TEMPR14[21] ), .D(sel_R_DATA_TEMPR15[21] ), .Y(
        OR4_131_Y));
    OR4 OR4_584 (.A(OR4_795_Y), .B(OR4_1022_Y), .C(OR4_597_Y), .D(
        OR4_386_Y), .Y(OR4_584_Y));
    OR4 OR4_659 (.A(sel_R_DATA_TEMPR20[22] ), .B(sel_R_DATA_TEMPR21[22] ), 
        .C(sel_R_DATA_TEMPR22[22] ), .D(sel_R_DATA_TEMPR23[22] ), .Y(
        OR4_659_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%3%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R3C0 (.A_DOUT({
        nc816, nc817, nc818, nc819, nc820,int_R_DATA_TEMPR3[31] , 
       int_R_DATA_TEMPR3[30] ,int_R_DATA_TEMPR3[29] ,int_R_DATA_TEMPR3[28] , 
       int_R_DATA_TEMPR3[27] ,int_R_DATA_TEMPR3[26] ,int_R_DATA_TEMPR3[25] , 
       int_R_DATA_TEMPR3[24] ,int_R_DATA_TEMPR3[23] ,int_R_DATA_TEMPR3[22] , 
       int_R_DATA_TEMPR3[21] ,int_R_DATA_TEMPR3[20] ,int_R_DATA_TEMPR3[19] , 
       int_R_DATA_TEMPR3[18] ,int_R_DATA_TEMPR3[17] }), .B_DOUT({nc821, 
        nc822, nc823,int_R_DATA_TEMPR3[16] ,int_R_DATA_TEMPR3[15] , 
       int_R_DATA_TEMPR3[14] ,int_R_DATA_TEMPR3[13] ,int_R_DATA_TEMPR3[12] , 
       int_R_DATA_TEMPR3[11] ,int_R_DATA_TEMPR3[10] ,int_R_DATA_TEMPR3[9] , 
       int_R_DATA_TEMPR3[8] ,int_R_DATA_TEMPR3[7] ,int_R_DATA_TEMPR3[6] , 
       int_R_DATA_TEMPR3[5] ,int_R_DATA_TEMPR3[4] ,int_R_DATA_TEMPR3[3] , 
       int_R_DATA_TEMPR3[2] ,int_R_DATA_TEMPR3[1] ,int_R_DATA_TEMPR3[0] }), 
        .DB_DETECT(int_DB_DETECT_NG[3] ), .SB_CORRECT( int_SB_CORRECT_NG[3] ), .ACCESS_BUSY(\ACCESS_BUSY[3] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[0] , R_ADDR[10], R_ADDR[9]}), .A_CLK(
        CLK), .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[0] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_982 (.A(sel_R_DATA_TEMPR96[13] ), .B(sel_R_DATA_TEMPR97[13] ), 
        .C(sel_R_DATA_TEMPR98[13] ), .D(sel_R_DATA_TEMPR99[13] ), .Y(
        OR4_982_Y));
    AND4 \AND4SB_CORRECT[72]  (.A(sel_SB_CORRECT_NG[72] ), .B(
        \BLKY2_pipe[18] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[72] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%13%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R13C0 (.A_DOUT({
        nc824, nc825, nc826, nc827, nc828,int_R_DATA_TEMPR13[31] , 
       int_R_DATA_TEMPR13[30] ,int_R_DATA_TEMPR13[29] , 
       int_R_DATA_TEMPR13[28] ,int_R_DATA_TEMPR13[27] , 
       int_R_DATA_TEMPR13[26] ,int_R_DATA_TEMPR13[25] , 
       int_R_DATA_TEMPR13[24] ,int_R_DATA_TEMPR13[23] , 
       int_R_DATA_TEMPR13[22] ,int_R_DATA_TEMPR13[21] , 
       int_R_DATA_TEMPR13[20] ,int_R_DATA_TEMPR13[19] , 
       int_R_DATA_TEMPR13[18] ,int_R_DATA_TEMPR13[17] }), .B_DOUT({nc829, 
        nc830, nc831,int_R_DATA_TEMPR13[16] ,int_R_DATA_TEMPR13[15] , 
       int_R_DATA_TEMPR13[14] ,int_R_DATA_TEMPR13[13] , 
       int_R_DATA_TEMPR13[12] ,int_R_DATA_TEMPR13[11] , 
       int_R_DATA_TEMPR13[10] ,int_R_DATA_TEMPR13[9] ,int_R_DATA_TEMPR13[8] , 
       int_R_DATA_TEMPR13[7] ,int_R_DATA_TEMPR13[6] ,int_R_DATA_TEMPR13[5] , 
       int_R_DATA_TEMPR13[4] ,int_R_DATA_TEMPR13[3] ,int_R_DATA_TEMPR13[2] , 
       int_R_DATA_TEMPR13[1] ,int_R_DATA_TEMPR13[0] }), .DB_DETECT( int_DB_DETECT_NG[13] ), .SB_CORRECT(int_SB_CORRECT_NG[13] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[13] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[3] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[3] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_596 (.A(sel_R_DATA_TEMPR112[28] ), .B(sel_R_DATA_TEMPR113[28] ), 
        .C(sel_R_DATA_TEMPR114[28] ), .D(sel_R_DATA_TEMPR115[28] ), .Y(
        OR4_596_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[8]  (.A(CFG3_13_Y), .B(CFG3_4_Y)
        , .Y(\BLKX2[8] ));
    OR4 OR4_256 (.A(OR4_994_Y), .B(OR4_880_Y), .C(OR4_816_Y), .D(
        OR4_296_Y), .Y(OR4_256_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%96%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R96C0 (.A_DOUT({
        nc832, nc833, nc834, nc835, nc836,int_R_DATA_TEMPR96[31] , 
       int_R_DATA_TEMPR96[30] ,int_R_DATA_TEMPR96[29] , 
       int_R_DATA_TEMPR96[28] ,int_R_DATA_TEMPR96[27] , 
       int_R_DATA_TEMPR96[26] ,int_R_DATA_TEMPR96[25] , 
       int_R_DATA_TEMPR96[24] ,int_R_DATA_TEMPR96[23] , 
       int_R_DATA_TEMPR96[22] ,int_R_DATA_TEMPR96[21] , 
       int_R_DATA_TEMPR96[20] ,int_R_DATA_TEMPR96[19] , 
       int_R_DATA_TEMPR96[18] ,int_R_DATA_TEMPR96[17] }), .B_DOUT({nc837, 
        nc838, nc839,int_R_DATA_TEMPR96[16] ,int_R_DATA_TEMPR96[15] , 
       int_R_DATA_TEMPR96[14] ,int_R_DATA_TEMPR96[13] , 
       int_R_DATA_TEMPR96[12] ,int_R_DATA_TEMPR96[11] , 
       int_R_DATA_TEMPR96[10] ,int_R_DATA_TEMPR96[9] ,int_R_DATA_TEMPR96[8] , 
       int_R_DATA_TEMPR96[7] ,int_R_DATA_TEMPR96[6] ,int_R_DATA_TEMPR96[5] , 
       int_R_DATA_TEMPR96[4] ,int_R_DATA_TEMPR96[3] ,int_R_DATA_TEMPR96[2] , 
       int_R_DATA_TEMPR96[1] ,int_R_DATA_TEMPR96[0] }), .DB_DETECT( int_DB_DETECT_NG[96] ), .SB_CORRECT(int_SB_CORRECT_NG[96] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[96] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[24] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[24] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR2 OR2_0 (.A(sel_R_DATA_TEMPR84[16] ), .B(sel_R_DATA_TEMPR85[16] ), .Y(
        OR2_0_Y));
    OR4 OR4_1255 (.A(sel_R_DATA_TEMPR12[14] ), .B(sel_R_DATA_TEMPR13[14] ), 
        .C(sel_R_DATA_TEMPR14[14] ), .D(sel_R_DATA_TEMPR15[14] ), .Y(
        OR4_1255_Y));
    AND4 \AND4DB_DETECT[116]  (.A(sel_DB_DETECT_NG[116] ), .B(
        \BLKY2_pipe[29] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[116] ));
    OR4 OR4_1084 (.A(sel_R_DATA_TEMPR20[4] ), .B(sel_R_DATA_TEMPR21[4] ), .C(sel_R_DATA_TEMPR22[4] ), .D(sel_R_DATA_TEMPR23[4] ), .Y(OR4_1084_Y));
    OR4 OR4_75 (.A(sel_R_DATA_TEMPR108[12] ), .B(sel_R_DATA_TEMPR109[12] ), 
        .C(sel_R_DATA_TEMPR110[12] ), .D(sel_R_DATA_TEMPR111[12] ), .Y(
        OR4_75_Y));
    OR4 OR4_1248 (.A(sel_R_DATA_TEMPR8[29] ), .B(sel_R_DATA_TEMPR9[29] ), .C(sel_R_DATA_TEMPR10[29] ), .D(sel_R_DATA_TEMPR11[29] ), .Y(OR4_1248_Y)
        );
    OR2 OR2_6 (.A(sel_R_DATA_TEMPR84[28] ), .B(sel_R_DATA_TEMPR85[28] ), .Y(
        OR2_6_Y));
    OR4 OR4_1339 (.A(sel_R_DATA_TEMPR124[14] ), .B(sel_R_DATA_TEMPR125[14] ), 
        .C(sel_R_DATA_TEMPR126[14] ), .D(sel_R_DATA_TEMPR127[14] ), .Y(
        OR4_1339_Y));
    OR4 OR4_1263 (.A(OR4_1080_Y), .B(OR4_937_Y), .C(OR4_656_Y), .D(
        OR4_1070_Y), .Y(OR4_1263_Y));
    OR4 OR4_1227 (.A(sel_R_DATA_TEMPR68[7] ), .B(sel_R_DATA_TEMPR69[7] ), .C(sel_R_DATA_TEMPR70[7] ), .D(sel_R_DATA_TEMPR71[7] ), .Y(OR4_1227_Y));
    OR4 OR4_431 (.A(sel_R_DATA_TEMPR32[5] ), .B(sel_R_DATA_TEMPR33[5] ), .C(sel_R_DATA_TEMPR34[5] ), .D(sel_R_DATA_TEMPR35[5] ), .Y(OR4_431_Y));
    OR4 OR4_91 (.A(sel_R_DATA_TEMPR68[25] ), .B(sel_R_DATA_TEMPR69[25] ), .C(sel_R_DATA_TEMPR70[25] ), .D(sel_R_DATA_TEMPR71[25] ), .Y(OR4_91_Y));
    AND4 \AND4DB_DETECT[58]  (.A(sel_DB_DETECT_NG[58] ), .B(
        \BLKY2_pipe[14] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[58] ));
    CFG3 #( .INIT(8'h2) )  CFG3_2 (.A(R_EN), .B(R_ADDR[15]), .C(
        R_ADDR[14]), .Y(CFG3_2_Y));
    OR4 OR4_124 (.A(sel_R_DATA_TEMPR36[15] ), .B(sel_R_DATA_TEMPR37[15] ), 
        .C(sel_R_DATA_TEMPR38[15] ), .D(sel_R_DATA_TEMPR39[15] ), .Y(
        OR4_124_Y));
    OR4 OR4_438 (.A(sel_R_DATA_TEMPR68[13] ), .B(sel_R_DATA_TEMPR69[13] ), 
        .C(sel_R_DATA_TEMPR70[13] ), .D(sel_R_DATA_TEMPR71[13] ), .Y(
        OR4_438_Y));
    OR4 OR4_1383 (.A(sel_R_DATA_TEMPR100[7] ), .B(sel_R_DATA_TEMPR101[7] ), 
        .C(sel_R_DATA_TEMPR102[7] ), .D(sel_R_DATA_TEMPR103[7] ), .Y(
        OR4_1383_Y));
    OR4 OR4_1030 (.A(sel_R_DATA_TEMPR96[28] ), .B(sel_R_DATA_TEMPR97[28] ), 
        .C(sel_R_DATA_TEMPR98[28] ), .D(sel_R_DATA_TEMPR99[28] ), .Y(
        OR4_1030_Y));
    OR4 OR4_709 (.A(sel_R_DATA_TEMPR120[5] ), .B(sel_R_DATA_TEMPR121[5] ), 
        .C(sel_R_DATA_TEMPR122[5] ), .D(sel_R_DATA_TEMPR123[5] ), .Y(
        OR4_709_Y));
    OR4 OR4_381 (.A(sel_R_DATA_TEMPR24[4] ), .B(sel_R_DATA_TEMPR25[4] ), .C(sel_R_DATA_TEMPR26[4] ), .D(sel_R_DATA_TEMPR27[4] ), .Y(OR4_381_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[13]  (.D(\BLKY2[13] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[13] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%28%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R28C0 (.A_DOUT({
        nc840, nc841, nc842, nc843, nc844,int_R_DATA_TEMPR28[31] , 
       int_R_DATA_TEMPR28[30] ,int_R_DATA_TEMPR28[29] , 
       int_R_DATA_TEMPR28[28] ,int_R_DATA_TEMPR28[27] , 
       int_R_DATA_TEMPR28[26] ,int_R_DATA_TEMPR28[25] , 
       int_R_DATA_TEMPR28[24] ,int_R_DATA_TEMPR28[23] , 
       int_R_DATA_TEMPR28[22] ,int_R_DATA_TEMPR28[21] , 
       int_R_DATA_TEMPR28[20] ,int_R_DATA_TEMPR28[19] , 
       int_R_DATA_TEMPR28[18] ,int_R_DATA_TEMPR28[17] }), .B_DOUT({nc845, 
        nc846, nc847,int_R_DATA_TEMPR28[16] ,int_R_DATA_TEMPR28[15] , 
       int_R_DATA_TEMPR28[14] ,int_R_DATA_TEMPR28[13] , 
       int_R_DATA_TEMPR28[12] ,int_R_DATA_TEMPR28[11] , 
       int_R_DATA_TEMPR28[10] ,int_R_DATA_TEMPR28[9] ,int_R_DATA_TEMPR28[8] , 
       int_R_DATA_TEMPR28[7] ,int_R_DATA_TEMPR28[6] ,int_R_DATA_TEMPR28[5] , 
       int_R_DATA_TEMPR28[4] ,int_R_DATA_TEMPR28[3] ,int_R_DATA_TEMPR28[2] , 
       int_R_DATA_TEMPR28[1] ,int_R_DATA_TEMPR28[0] }), .DB_DETECT( int_DB_DETECT_NG[28] ), .SB_CORRECT(int_SB_CORRECT_NG[28] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[28] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[7] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[24]  (.A(CFG3_16_Y), .B(
        CFG3_3_Y), .Y(\BLKY2[24] ));
    OR2 OR2_3 (.A(sel_R_DATA_TEMPR84[13] ), .B(sel_R_DATA_TEMPR85[13] ), .Y(
        OR2_3_Y));
    OR4 OR4_654 (.A(sel_R_DATA_TEMPR88[31] ), .B(sel_R_DATA_TEMPR89[31] ), 
        .C(sel_R_DATA_TEMPR90[31] ), .D(sel_R_DATA_TEMPR91[31] ), .Y(
        OR4_654_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%25%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R25C0 (.A_DOUT({
        nc848, nc849, nc850, nc851, nc852,int_R_DATA_TEMPR25[31] , 
       int_R_DATA_TEMPR25[30] ,int_R_DATA_TEMPR25[29] , 
       int_R_DATA_TEMPR25[28] ,int_R_DATA_TEMPR25[27] , 
       int_R_DATA_TEMPR25[26] ,int_R_DATA_TEMPR25[25] , 
       int_R_DATA_TEMPR25[24] ,int_R_DATA_TEMPR25[23] , 
       int_R_DATA_TEMPR25[22] ,int_R_DATA_TEMPR25[21] , 
       int_R_DATA_TEMPR25[20] ,int_R_DATA_TEMPR25[19] , 
       int_R_DATA_TEMPR25[18] ,int_R_DATA_TEMPR25[17] }), .B_DOUT({nc853, 
        nc854, nc855,int_R_DATA_TEMPR25[16] ,int_R_DATA_TEMPR25[15] , 
       int_R_DATA_TEMPR25[14] ,int_R_DATA_TEMPR25[13] , 
       int_R_DATA_TEMPR25[12] ,int_R_DATA_TEMPR25[11] , 
       int_R_DATA_TEMPR25[10] ,int_R_DATA_TEMPR25[9] ,int_R_DATA_TEMPR25[8] , 
       int_R_DATA_TEMPR25[7] ,int_R_DATA_TEMPR25[6] ,int_R_DATA_TEMPR25[5] , 
       int_R_DATA_TEMPR25[4] ,int_R_DATA_TEMPR25[3] ,int_R_DATA_TEMPR25[2] , 
       int_R_DATA_TEMPR25[1] ,int_R_DATA_TEMPR25[0] }), .DB_DETECT( int_DB_DETECT_NG[25] ), .SB_CORRECT(int_SB_CORRECT_NG[25] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[25] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[6] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_947 (.A(sel_R_DATA_TEMPR120[13] ), .B(sel_R_DATA_TEMPR121[13] ), 
        .C(sel_R_DATA_TEMPR122[13] ), .D(sel_R_DATA_TEMPR123[13] ), .Y(
        OR4_947_Y));
    OR4 OR4_804 (.A(sel_R_DATA_TEMPR80[30] ), .B(sel_R_DATA_TEMPR81[30] ), 
        .C(sel_R_DATA_TEMPR82[30] ), .D(sel_R_DATA_TEMPR83[30] ), .Y(
        OR4_804_Y));
    OR4 OR4_779 (.A(OR4_583_Y), .B(OR4_320_Y), .C(OR4_672_Y), .D(
        OR4_528_Y), .Y(OR4_779_Y));
    OR4 OR4_1324 (.A(sel_R_DATA_TEMPR116[18] ), .B(sel_R_DATA_TEMPR117[18] ), 
        .C(sel_R_DATA_TEMPR118[18] ), .D(sel_R_DATA_TEMPR119[18] ), .Y(
        OR4_1324_Y));
    OR4 OR4_923 (.A(sel_R_DATA_TEMPR40[4] ), .B(sel_R_DATA_TEMPR41[4] ), .C(sel_R_DATA_TEMPR42[4] ), .D(sel_R_DATA_TEMPR43[4] ), .Y(OR4_923_Y));
    OR4 OR4_480 (.A(sel_R_DATA_TEMPR36[4] ), .B(sel_R_DATA_TEMPR37[4] ), .C(sel_R_DATA_TEMPR38[4] ), .D(sel_R_DATA_TEMPR39[4] ), .Y(OR4_480_Y));
    OR4 OR4_503 (.A(OR4_87_Y), .B(OR4_344_Y), .C(OR4_547_Y), .D(
        OR4_387_Y), .Y(OR4_503_Y));
    OR4 OR4_314 (.A(sel_R_DATA_TEMPR16[24] ), .B(sel_R_DATA_TEMPR17[24] ), 
        .C(sel_R_DATA_TEMPR18[24] ), .D(sel_R_DATA_TEMPR19[24] ), .Y(
        OR4_314_Y));
    CFG3 #( .INIT(8'h80) )  CFG3_21 (.A(R_ADDR[13]), .B(R_ADDR[12]), 
        .C(R_ADDR[11]), .Y(CFG3_21_Y));
    OR4 OR4_1006 (.A(sel_R_DATA_TEMPR44[24] ), .B(sel_R_DATA_TEMPR45[24] ), 
        .C(sel_R_DATA_TEMPR46[24] ), .D(sel_R_DATA_TEMPR47[24] ), .Y(
        OR4_1006_Y));
    OR4 OR4_874 (.A(sel_R_DATA_TEMPR76[13] ), .B(sel_R_DATA_TEMPR77[13] ), 
        .C(sel_R_DATA_TEMPR78[13] ), .D(sel_R_DATA_TEMPR79[13] ), .Y(
        OR4_874_Y));
    OR4 OR4_826 (.A(sel_R_DATA_TEMPR48[10] ), .B(sel_R_DATA_TEMPR49[10] ), 
        .C(sel_R_DATA_TEMPR50[10] ), .D(sel_R_DATA_TEMPR51[10] ), .Y(
        OR4_826_Y));
    OR4 OR4_721 (.A(sel_R_DATA_TEMPR80[6] ), .B(sel_R_DATA_TEMPR81[6] ), .C(sel_R_DATA_TEMPR82[6] ), .D(sel_R_DATA_TEMPR83[6] ), .Y(OR4_721_Y));
    OR4 OR4_43 (.A(sel_R_DATA_TEMPR24[31] ), .B(sel_R_DATA_TEMPR25[31] ), .C(sel_R_DATA_TEMPR26[31] ), .D(sel_R_DATA_TEMPR27[31] ), .Y(OR4_43_Y));
    OR4 OR4_1169 (.A(sel_R_DATA_TEMPR48[15] ), .B(sel_R_DATA_TEMPR49[15] ), 
        .C(sel_R_DATA_TEMPR50[15] ), .D(sel_R_DATA_TEMPR51[15] ), .Y(
        OR4_1169_Y));
    OR4 OR4_573 (.A(sel_R_DATA_TEMPR112[19] ), .B(sel_R_DATA_TEMPR113[19] ), 
        .C(sel_R_DATA_TEMPR114[19] ), .D(sel_R_DATA_TEMPR115[19] ), .Y(
        OR4_573_Y));
    OR4 OR4_539 (.A(sel_R_DATA_TEMPR56[17] ), .B(sel_R_DATA_TEMPR57[17] ), 
        .C(sel_R_DATA_TEMPR58[17] ), .D(sel_R_DATA_TEMPR59[17] ), .Y(
        OR4_539_Y));
    INV \INVBLKX0[0]  (.A(W_ADDR[9]), .Y(\BLKX0[0] ));
    OR2 OR2_26 (.A(sel_R_DATA_TEMPR84[20] ), .B(sel_R_DATA_TEMPR85[20] ), .Y(
        OR2_26_Y));
    OR4 OR4_111 (.A(OR4_1106_Y), .B(OR4_863_Y), .C(OR4_632_Y), .D(
        OR4_1337_Y), .Y(OR4_111_Y));
    OR4 OR4_598 (.A(OR4_363_Y), .B(OR4_201_Y), .C(OR4_1282_Y), .D(
        OR4_1135_Y), .Y(OR4_598_Y));
    CFG3 #( .INIT(8'h8) )  CFG3_1 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_1_Y));
    AND4 \AND4DB_DETECT[121]  (.A(sel_DB_DETECT_NG[121] ), .B(
        \BLKY2_pipe[30] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[121] ));
    AND4 \AND4DB_DETECT[75]  (.A(sel_DB_DETECT_NG[75] ), .B(
        \BLKY2_pipe[18] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[75] ));
    OR4 OR4_59 (.A(OR4_174_Y), .B(OR4_1202_Y), .C(OR4_917_Y), .D(
        OR4_1335_Y), .Y(OR4_59_Y));
    AND4 \AND4SB_CORRECT[111]  (.A(sel_SB_CORRECT_NG[111] ), .B(
        \BLKY2_pipe[27] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[111] ));
    OR4 OR4_530 (.A(sel_R_DATA_TEMPR52[14] ), .B(sel_R_DATA_TEMPR53[14] ), 
        .C(sel_R_DATA_TEMPR54[14] ), .D(sel_R_DATA_TEMPR55[14] ), .Y(
        OR4_530_Y));
    OR4 OR4_1301 (.A(sel_R_DATA_TEMPR120[7] ), .B(sel_R_DATA_TEMPR121[7] ), 
        .C(sel_R_DATA_TEMPR122[7] ), .D(sel_R_DATA_TEMPR123[7] ), .Y(
        OR4_1301_Y));
    AND4 \AND4SB_CORRECT[52]  (.A(sel_SB_CORRECT_NG[52] ), .B(
        \BLKY2_pipe[13] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[52] ));
    OR4 OR4_263 (.A(OR4_244_Y), .B(OR2_19_Y), .C(sel_R_DATA_TEMPR86[5] ), 
        .D(sel_R_DATA_TEMPR87[5] ), .Y(OR4_263_Y));
    OR4 OR4_526 (.A(\SB_CORRECT[104] ), .B(\SB_CORRECT[105] ), 
        .C(\SB_CORRECT[106] ), .D(\SB_CORRECT[107] ), .Y(
        OR4_526_Y));
    OR4 OR4_1293 (.A(sel_R_DATA_TEMPR8[6] ), .B(sel_R_DATA_TEMPR9[6] ), .C(sel_R_DATA_TEMPR10[6] ), .D(sel_R_DATA_TEMPR11[6] ), .Y(OR4_1293_Y));
    OR4 OR4_1145 (.A(sel_R_DATA_TEMPR108[6] ), .B(sel_R_DATA_TEMPR109[6] ), 
        .C(sel_R_DATA_TEMPR110[6] ), .D(sel_R_DATA_TEMPR111[6] ), .Y(
        OR4_1145_Y));
    AND4 \AND4SB_CORRECT[30]  (.A(sel_SB_CORRECT_NG[30] ), .B(
        \BLKY2_pipe[7] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[30] ));
    OR4 OR4_445 (.A(sel_R_DATA_TEMPR124[11] ), .B(sel_R_DATA_TEMPR125[11] ), 
        .C(sel_R_DATA_TEMPR126[11] ), .D(sel_R_DATA_TEMPR127[11] ), .Y(
        OR4_445_Y));
    OR4 OR4_1329 (.A(sel_R_DATA_TEMPR28[11] ), .B(sel_R_DATA_TEMPR29[11] ), 
        .C(sel_R_DATA_TEMPR30[11] ), .D(sel_R_DATA_TEMPR31[11] ), .Y(
        OR4_1329_Y));
    OR4 OR4_411 (.A(sel_R_DATA_TEMPR88[14] ), .B(sel_R_DATA_TEMPR89[14] ), 
        .C(sel_R_DATA_TEMPR90[14] ), .D(sel_R_DATA_TEMPR91[14] ), .Y(
        OR4_411_Y));
    OR4 OR4_1041 (.A(OR4_142_Y), .B(OR4_580_Y), .C(OR4_170_Y), .D(
        OR4_1130_Y), .Y(OR4_1041_Y));
    CFG3 #( .INIT(8'h20) )  CFG3_11 (.A(R_ADDR[13]), .B(R_ADDR[12]), 
        .C(R_ADDR[11]), .Y(CFG3_11_Y));
    OR4 OR4_496 (.A(OR4_609_Y), .B(OR4_828_Y), .C(OR4_426_Y), .D(
        OR4_198_Y), .Y(OR4_496_Y));
    OR4 OR4_418 (.A(OR4_362_Y), .B(OR4_1084_Y), .C(OR4_381_Y), .D(
        OR4_590_Y), .Y(OR4_418_Y));
    OR4 OR4_1086 (.A(OR4_254_Y), .B(OR4_1047_Y), .C(OR4_1116_Y), .D(
        OR4_436_Y), .Y(OR4_1086_Y));
    OR4 OR4_1020 (.A(OR4_533_Y), .B(OR4_1210_Y), .C(OR4_208_Y), .D(
        OR4_477_Y), .Y(OR4_1020_Y));
    AND4 \AND4SB_CORRECT[117]  (.A(sel_SB_CORRECT_NG[117] ), .B(
        \BLKY2_pipe[29] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[117] ));
    OR4 OR4_968 (.A(sel_R_DATA_TEMPR8[14] ), .B(sel_R_DATA_TEMPR9[14] ), .C(sel_R_DATA_TEMPR10[14] ), .D(sel_R_DATA_TEMPR11[14] ), .Y(OR4_968_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%41%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R41C0 (.A_DOUT({
        nc856, nc857, nc858, nc859, nc860,int_R_DATA_TEMPR41[31] , 
       int_R_DATA_TEMPR41[30] ,int_R_DATA_TEMPR41[29] , 
       int_R_DATA_TEMPR41[28] ,int_R_DATA_TEMPR41[27] , 
       int_R_DATA_TEMPR41[26] ,int_R_DATA_TEMPR41[25] , 
       int_R_DATA_TEMPR41[24] ,int_R_DATA_TEMPR41[23] , 
       int_R_DATA_TEMPR41[22] ,int_R_DATA_TEMPR41[21] , 
       int_R_DATA_TEMPR41[20] ,int_R_DATA_TEMPR41[19] , 
       int_R_DATA_TEMPR41[18] ,int_R_DATA_TEMPR41[17] }), .B_DOUT({nc861, 
        nc862, nc863,int_R_DATA_TEMPR41[16] ,int_R_DATA_TEMPR41[15] , 
       int_R_DATA_TEMPR41[14] ,int_R_DATA_TEMPR41[13] , 
       int_R_DATA_TEMPR41[12] ,int_R_DATA_TEMPR41[11] , 
       int_R_DATA_TEMPR41[10] ,int_R_DATA_TEMPR41[9] ,int_R_DATA_TEMPR41[8] , 
       int_R_DATA_TEMPR41[7] ,int_R_DATA_TEMPR41[6] ,int_R_DATA_TEMPR41[5] , 
       int_R_DATA_TEMPR41[4] ,int_R_DATA_TEMPR41[3] ,int_R_DATA_TEMPR41[2] , 
       int_R_DATA_TEMPR41[1] ,int_R_DATA_TEMPR41[0] }), .DB_DETECT( int_DB_DETECT_NG[41] ), .SB_CORRECT(int_SB_CORRECT_NG[41] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[41] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[10] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[10] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4DB_DETECT[123]  (.A(sel_DB_DETECT_NG[123] ), .B(
        \BLKY2_pipe[30] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[123] ));
    DFN1E1 \DFN1E1BLKY2_pipe[12]  (.D(\BLKY2[12] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[12] ));
    OR4 OR4_1166 (.A(OR4_276_Y), .B(OR4_530_Y), .C(OR4_732_Y), .D(
        OR4_568_Y), .Y(OR4_1166_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%50%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R50C0 (.A_DOUT({
        nc864, nc865, nc866, nc867, nc868,int_R_DATA_TEMPR50[31] , 
       int_R_DATA_TEMPR50[30] ,int_R_DATA_TEMPR50[29] , 
       int_R_DATA_TEMPR50[28] ,int_R_DATA_TEMPR50[27] , 
       int_R_DATA_TEMPR50[26] ,int_R_DATA_TEMPR50[25] , 
       int_R_DATA_TEMPR50[24] ,int_R_DATA_TEMPR50[23] , 
       int_R_DATA_TEMPR50[22] ,int_R_DATA_TEMPR50[21] , 
       int_R_DATA_TEMPR50[20] ,int_R_DATA_TEMPR50[19] , 
       int_R_DATA_TEMPR50[18] ,int_R_DATA_TEMPR50[17] }), .B_DOUT({nc869, 
        nc870, nc871,int_R_DATA_TEMPR50[16] ,int_R_DATA_TEMPR50[15] , 
       int_R_DATA_TEMPR50[14] ,int_R_DATA_TEMPR50[13] , 
       int_R_DATA_TEMPR50[12] ,int_R_DATA_TEMPR50[11] , 
       int_R_DATA_TEMPR50[10] ,int_R_DATA_TEMPR50[9] ,int_R_DATA_TEMPR50[8] , 
       int_R_DATA_TEMPR50[7] ,int_R_DATA_TEMPR50[6] ,int_R_DATA_TEMPR50[5] , 
       int_R_DATA_TEMPR50[4] ,int_R_DATA_TEMPR50[3] ,int_R_DATA_TEMPR50[2] , 
       int_R_DATA_TEMPR50[1] ,int_R_DATA_TEMPR50[0] }), .DB_DETECT( int_DB_DETECT_NG[50] ), .SB_CORRECT(int_SB_CORRECT_NG[50] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[50] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[12] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[12] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1381 (.A(sel_R_DATA_TEMPR12[12] ), .B(sel_R_DATA_TEMPR13[12] ), 
        .C(sel_R_DATA_TEMPR14[12] ), .D(sel_R_DATA_TEMPR15[12] ), .Y(
        OR4_1381_Y));
    OR4 \OR4_R_DATA[0]  (.A(OR4_1142_Y), .B(OR4_1305_Y), .C(OR4_854_Y), 
        .D(OR4_1129_Y), .Y(R_DATA[0]));
    OR4 OR4_389 (.A(sel_R_DATA_TEMPR20[11] ), .B(sel_R_DATA_TEMPR21[11] ), 
        .C(sel_R_DATA_TEMPR22[11] ), .D(sel_R_DATA_TEMPR23[11] ), .Y(
        OR4_389_Y));
    OR4 OR4_1261 (.A(sel_R_DATA_TEMPR12[2] ), .B(sel_R_DATA_TEMPR13[2] ), .C(sel_R_DATA_TEMPR14[2] ), .D(sel_R_DATA_TEMPR15[2] ), .Y(OR4_1261_Y));
    OR4 OR4_392 (.A(\DB_DETECT[64] ), .B(\DB_DETECT[65] ), .C(
        \DB_DETECT[66] ), .D(\DB_DETECT[67] ), .Y(OR4_392_Y));
    OR4 OR4_1043 (.A(sel_R_DATA_TEMPR60[21] ), .B(sel_R_DATA_TEMPR61[21] ), 
        .C(sel_R_DATA_TEMPR62[21] ), .D(sel_R_DATA_TEMPR63[21] ), .Y(
        OR4_1043_Y));
    OR4 OR4_1168 (.A(sel_R_DATA_TEMPR104[27] ), .B(sel_R_DATA_TEMPR105[27] ), 
        .C(sel_R_DATA_TEMPR106[27] ), .D(sel_R_DATA_TEMPR107[27] ), .Y(
        OR4_1168_Y));
    OR4 OR4_1199 (.A(sel_R_DATA_TEMPR92[6] ), .B(sel_R_DATA_TEMPR93[6] ), .C(sel_R_DATA_TEMPR94[6] ), .D(sel_R_DATA_TEMPR95[6] ), .Y(OR4_1199_Y));
    OR4 OR4_19 (.A(sel_R_DATA_TEMPR28[27] ), .B(sel_R_DATA_TEMPR29[27] ), .C(sel_R_DATA_TEMPR30[27] ), .D(sel_R_DATA_TEMPR31[27] ), .Y(OR4_19_Y));
    OR4 OR4_41 (.A(sel_R_DATA_TEMPR68[19] ), .B(sel_R_DATA_TEMPR69[19] ), .C(sel_R_DATA_TEMPR70[19] ), .D(sel_R_DATA_TEMPR71[19] ), .Y(OR4_41_Y));
    OR4 OR4_333 (.A(OR4_98_Y), .B(OR4_86_Y), .C(OR4_527_Y), .D(
        OR4_916_Y), .Y(OR4_333_Y));
    OR4 OR4_730 (.A(sel_R_DATA_TEMPR124[30] ), .B(sel_R_DATA_TEMPR125[30] ), 
        .C(sel_R_DATA_TEMPR126[30] ), .D(sel_R_DATA_TEMPR127[30] ), .Y(
        OR4_730_Y));
    OR4 OR4_519 (.A(sel_R_DATA_TEMPR124[27] ), .B(sel_R_DATA_TEMPR125[27] ), 
        .C(sel_R_DATA_TEMPR126[27] ), .D(sel_R_DATA_TEMPR127[27] ), .Y(
        OR4_519_Y));
    OR4 OR4_1279 (.A(OR4_357_Y), .B(OR4_584_Y), .C(OR4_578_Y), .D(
        OR4_806_Y), .Y(OR4_1279_Y));
    OR4 OR4_668 (.A(sel_R_DATA_TEMPR112[21] ), .B(sel_R_DATA_TEMPR113[21] ), 
        .C(sel_R_DATA_TEMPR114[21] ), .D(sel_R_DATA_TEMPR115[21] ), .Y(
        OR4_668_Y));
    OR4 OR4_510 (.A(OR4_495_Y), .B(OR4_275_Y), .C(OR4_24_Y), .D(
        OR4_39_Y), .Y(OR4_510_Y));
    AND4 \AND4DB_DETECT[88]  (.A(sel_DB_DETECT_NG[88] ), .B(
        \BLKY2_pipe[22] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[88] ));
    OR4 OR4_1054 (.A(sel_R_DATA_TEMPR48[21] ), .B(sel_R_DATA_TEMPR49[21] ), 
        .C(sel_R_DATA_TEMPR50[21] ), .D(sel_R_DATA_TEMPR51[21] ), .Y(
        OR4_1054_Y));
    OR4 OR4_444 (.A(sel_R_DATA_TEMPR104[15] ), .B(sel_R_DATA_TEMPR105[15] ), 
        .C(sel_R_DATA_TEMPR106[15] ), .D(sel_R_DATA_TEMPR107[15] ), .Y(
        OR4_444_Y));
    OR4 OR4_432 (.A(\SB_CORRECT[4] ), .B(\SB_CORRECT[5] ), .C(
        \SB_CORRECT[6] ), .D(\SB_CORRECT[7] ), .Y(OR4_432_Y));
    OR4 OR4_528 (.A(sel_R_DATA_TEMPR12[31] ), .B(sel_R_DATA_TEMPR13[31] ), 
        .C(sel_R_DATA_TEMPR14[31] ), .D(sel_R_DATA_TEMPR15[31] ), .Y(
        OR4_528_Y));
    AND4 \AND4DB_DETECT[59]  (.A(sel_DB_DETECT_NG[59] ), .B(
        \BLKY2_pipe[14] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[59] ));
    OR4 OR4_52 (.A(sel_R_DATA_TEMPR52[0] ), .B(sel_R_DATA_TEMPR53[0] ), .C(sel_R_DATA_TEMPR54[0] ), .D(sel_R_DATA_TEMPR55[0] ), .Y(OR4_52_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[2]  (.D(\BLKY2[2] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[2] ));
    OR4 OR4_1353 (.A(OR4_147_Y), .B(OR4_419_Y), .C(OR4_610_Y), .D(
        OR4_463_Y), .Y(OR4_1353_Y));
    OR4 OR4_1131 (.A(OR4_1020_Y), .B(OR4_722_Y), .C(OR4_1033_Y), .D(
        OR4_288_Y), .Y(OR4_1131_Y));
    OR4 OR4_662 (.A(sel_R_DATA_TEMPR88[9] ), .B(sel_R_DATA_TEMPR89[9] ), .C(sel_R_DATA_TEMPR90[9] ), .D(sel_R_DATA_TEMPR91[9] ), .Y(OR4_662_Y));
    OR4 OR4_439 (.A(OR4_1175_Y), .B(OR2_12_Y), .C(sel_R_DATA_TEMPR86[18] )
        , .D(sel_R_DATA_TEMPR87[18] ), .Y(OR4_439_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_18 (.A(R_ADDR[13]), .B(R_ADDR[12]), .C(
        R_ADDR[11]), .Y(CFG3_18_Y));
    OR4 OR4_346 (.A(sel_R_DATA_TEMPR12[11] ), .B(sel_R_DATA_TEMPR13[11] ), 
        .C(sel_R_DATA_TEMPR14[11] ), .D(sel_R_DATA_TEMPR15[11] ), .Y(
        OR4_346_Y));
    OR2 OR2_20 (.A(sel_R_DATA_TEMPR84[11] ), .B(sel_R_DATA_TEMPR85[11] ), .Y(
        OR2_20_Y));
    OR4 OR4_136 (.A(sel_R_DATA_TEMPR32[21] ), .B(sel_R_DATA_TEMPR33[21] ), 
        .C(sel_R_DATA_TEMPR34[21] ), .D(sel_R_DATA_TEMPR35[21] ), .Y(
        OR4_136_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%89%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R89C0 (.A_DOUT({
        nc872, nc873, nc874, nc875, nc876,int_R_DATA_TEMPR89[31] , 
       int_R_DATA_TEMPR89[30] ,int_R_DATA_TEMPR89[29] , 
       int_R_DATA_TEMPR89[28] ,int_R_DATA_TEMPR89[27] , 
       int_R_DATA_TEMPR89[26] ,int_R_DATA_TEMPR89[25] , 
       int_R_DATA_TEMPR89[24] ,int_R_DATA_TEMPR89[23] , 
       int_R_DATA_TEMPR89[22] ,int_R_DATA_TEMPR89[21] , 
       int_R_DATA_TEMPR89[20] ,int_R_DATA_TEMPR89[19] , 
       int_R_DATA_TEMPR89[18] ,int_R_DATA_TEMPR89[17] }), .B_DOUT({nc877, 
        nc878, nc879,int_R_DATA_TEMPR89[16] ,int_R_DATA_TEMPR89[15] , 
       int_R_DATA_TEMPR89[14] ,int_R_DATA_TEMPR89[13] , 
       int_R_DATA_TEMPR89[12] ,int_R_DATA_TEMPR89[11] , 
       int_R_DATA_TEMPR89[10] ,int_R_DATA_TEMPR89[9] ,int_R_DATA_TEMPR89[8] , 
       int_R_DATA_TEMPR89[7] ,int_R_DATA_TEMPR89[6] ,int_R_DATA_TEMPR89[5] , 
       int_R_DATA_TEMPR89[4] ,int_R_DATA_TEMPR89[3] ,int_R_DATA_TEMPR89[2] , 
       int_R_DATA_TEMPR89[1] ,int_R_DATA_TEMPR89[0] }), .DB_DETECT( int_DB_DETECT_NG[89] ), .SB_CORRECT(int_SB_CORRECT_NG[89] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[89] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[22] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[22] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1315 (.A(OR4_490_Y), .B(OR4_1151_Y), .C(OR4_153_Y), .D(
        OR4_428_Y), .Y(OR4_1315_Y));
    INV \INVBLKX1[0]  (.A(W_ADDR[10]), .Y(\BLKX1[0] ));
    DFN1E1 \DFN1E1BLKY2_pipe[6]  (.D(\BLKY2[6] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[6] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%62%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R62C0 (.A_DOUT({
        nc880, nc881, nc882, nc883, nc884,int_R_DATA_TEMPR62[31] , 
       int_R_DATA_TEMPR62[30] ,int_R_DATA_TEMPR62[29] , 
       int_R_DATA_TEMPR62[28] ,int_R_DATA_TEMPR62[27] , 
       int_R_DATA_TEMPR62[26] ,int_R_DATA_TEMPR62[25] , 
       int_R_DATA_TEMPR62[24] ,int_R_DATA_TEMPR62[23] , 
       int_R_DATA_TEMPR62[22] ,int_R_DATA_TEMPR62[21] , 
       int_R_DATA_TEMPR62[20] ,int_R_DATA_TEMPR62[19] , 
       int_R_DATA_TEMPR62[18] ,int_R_DATA_TEMPR62[17] }), .B_DOUT({nc885, 
        nc886, nc887,int_R_DATA_TEMPR62[16] ,int_R_DATA_TEMPR62[15] , 
       int_R_DATA_TEMPR62[14] ,int_R_DATA_TEMPR62[13] , 
       int_R_DATA_TEMPR62[12] ,int_R_DATA_TEMPR62[11] , 
       int_R_DATA_TEMPR62[10] ,int_R_DATA_TEMPR62[9] ,int_R_DATA_TEMPR62[8] , 
       int_R_DATA_TEMPR62[7] ,int_R_DATA_TEMPR62[6] ,int_R_DATA_TEMPR62[5] , 
       int_R_DATA_TEMPR62[4] ,int_R_DATA_TEMPR62[3] ,int_R_DATA_TEMPR62[2] , 
       int_R_DATA_TEMPR62[1] ,int_R_DATA_TEMPR62[0] }), .DB_DETECT( int_DB_DETECT_NG[62] ), .SB_CORRECT(int_SB_CORRECT_NG[62] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[62] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[15] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[15] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR2 OR2_16 (.A(sel_R_DATA_TEMPR84[30] ), .B(sel_R_DATA_TEMPR85[30] ), .Y(
        OR2_16_Y));
    CFG3 #( .INIT(8'h20) )  CFG3_22 (.A(W_ADDR[13]), .B(W_ADDR[12]), 
        .C(W_ADDR[11]), .Y(CFG3_22_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[20]  (.A(CFG3_18_Y), .B(
        CFG3_9_Y), .Y(\BLKY2[20] ));
    OR2 OR2_27 (.A(sel_R_DATA_TEMPR84[6] ), .B(sel_R_DATA_TEMPR85[6] ), .Y(
        OR2_27_Y));
    AND4 \AND4SB_CORRECT[43]  (.A(sel_SB_CORRECT_NG[43] ), .B(
        \BLKY2_pipe[10] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[43] ));
    OR4 OR4_426 (.A(sel_R_DATA_TEMPR24[28] ), .B(sel_R_DATA_TEMPR25[28] ), 
        .C(sel_R_DATA_TEMPR26[28] ), .D(sel_R_DATA_TEMPR27[28] ), .Y(
        OR4_426_Y));
    OR4 OR4_1196 (.A(sel_R_DATA_TEMPR28[8] ), .B(sel_R_DATA_TEMPR29[8] ), .C(sel_R_DATA_TEMPR30[8] ), .D(sel_R_DATA_TEMPR31[8] ), .Y(OR4_1196_Y));
    OR4 OR4_203 (.A(sel_R_DATA_TEMPR76[31] ), .B(sel_R_DATA_TEMPR77[31] ), 
        .C(sel_R_DATA_TEMPR78[31] ), .D(sel_R_DATA_TEMPR79[31] ), .Y(
        OR4_203_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[19]  (.A(CFG3_5_Y), .B(
        CFG3_17_Y), .Y(\BLKX2[19] ));
    OR4 OR4_290 (.A(sel_R_DATA_TEMPR104[9] ), .B(sel_R_DATA_TEMPR105[9] ), 
        .C(sel_R_DATA_TEMPR106[9] ), .D(sel_R_DATA_TEMPR107[9] ), .Y(
        OR4_290_Y));
    OR4 OR4_597 (.A(sel_R_DATA_TEMPR24[21] ), .B(sel_R_DATA_TEMPR25[21] ), 
        .C(sel_R_DATA_TEMPR26[21] ), .D(sel_R_DATA_TEMPR27[21] ), .Y(
        OR4_597_Y));
    AND4 \AND4DB_DETECT[6]  (.A(sel_DB_DETECT_NG[6] ), .B(
        \BLKY2_pipe[1] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[6] ));
    AND4 \AND4SB_CORRECT[4]  (.A(sel_SB_CORRECT_NG[4] ), .B(
        \BLKY2_pipe[1] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[4] ));
    OR4 OR4_1102 (.A(sel_R_DATA_TEMPR20[26] ), .B(sel_R_DATA_TEMPR21[26] ), 
        .C(sel_R_DATA_TEMPR22[26] ), .D(sel_R_DATA_TEMPR23[26] ), .Y(
        OR4_1102_Y));
    OR4 OR4_1291 (.A(sel_R_DATA_TEMPR52[30] ), .B(sel_R_DATA_TEMPR53[30] ), 
        .C(sel_R_DATA_TEMPR54[30] ), .D(sel_R_DATA_TEMPR55[30] ), .Y(
        OR4_1291_Y));
    OR4 OR4_858 (.A(sel_R_DATA_TEMPR56[16] ), .B(sel_R_DATA_TEMPR57[16] ), 
        .C(sel_R_DATA_TEMPR58[16] ), .D(sel_R_DATA_TEMPR59[16] ), .Y(
        OR4_858_Y));
    OR4 OR4_789 (.A(sel_R_DATA_TEMPR24[2] ), .B(sel_R_DATA_TEMPR25[2] ), .C(sel_R_DATA_TEMPR26[2] ), .D(sel_R_DATA_TEMPR27[2] ), .Y(OR4_789_Y));
    OR4 OR4_338 (.A(sel_R_DATA_TEMPR52[17] ), .B(sel_R_DATA_TEMPR53[17] ), 
        .C(sel_R_DATA_TEMPR54[17] ), .D(sel_R_DATA_TEMPR55[17] ), .Y(
        OR4_338_Y));
    OR4 OR4_273 (.A(sel_R_DATA_TEMPR32[20] ), .B(sel_R_DATA_TEMPR33[20] ), 
        .C(sel_R_DATA_TEMPR34[20] ), .D(sel_R_DATA_TEMPR35[20] ), .Y(
        OR4_273_Y));
    OR4 OR4_1198 (.A(OR4_505_Y), .B(OR4_1380_Y), .C(OR4_195_Y), .D(
        OR4_676_Y), .Y(OR4_1198_Y));
    OR4 OR4_908 (.A(sel_R_DATA_TEMPR48[12] ), .B(sel_R_DATA_TEMPR49[12] ), 
        .C(sel_R_DATA_TEMPR50[12] ), .D(sel_R_DATA_TEMPR51[12] ), .Y(
        OR4_908_Y));
    AND4 \AND4SB_CORRECT[95]  (.A(sel_SB_CORRECT_NG[95] ), .B(
        \BLKY2_pipe[23] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[95] ));
    AND4 \AND4SB_CORRECT[96]  (.A(sel_SB_CORRECT_NG[96] ), .B(
        \BLKY2_pipe[24] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[96] ));
    OR4 OR4_313 (.A(OR4_558_Y), .B(OR4_1044_Y), .C(OR4_334_Y), .D(
        OR4_548_Y), .Y(OR4_313_Y));
    OR4 OR4_322 (.A(sel_R_DATA_TEMPR100[0] ), .B(sel_R_DATA_TEMPR101[0] ), 
        .C(sel_R_DATA_TEMPR102[0] ), .D(sel_R_DATA_TEMPR103[0] ), .Y(
        OR4_322_Y));
    OR4 OR4_865 (.A(OR4_1275_Y), .B(OR4_1336_Y), .C(OR4_355_Y), .D(
        OR4_240_Y), .Y(OR4_865_Y));
    OR4 OR4_710 (.A(OR4_561_Y), .B(OR4_359_Y), .C(OR4_803_Y), .D(
        OR4_1205_Y), .Y(OR4_710_Y));
    OR4 OR4_1048 (.A(sel_R_DATA_TEMPR56[2] ), .B(sel_R_DATA_TEMPR57[2] ), .C(sel_R_DATA_TEMPR58[2] ), .D(sel_R_DATA_TEMPR59[2] ), .Y(OR4_1048_Y));
    OR4 OR4_884 (.A(sel_R_DATA_TEMPR12[13] ), .B(sel_R_DATA_TEMPR13[13] ), 
        .C(sel_R_DATA_TEMPR14[13] ), .D(sel_R_DATA_TEMPR15[13] ), .Y(
        OR4_884_Y));
    OR4 OR4_699 (.A(OR4_549_Y), .B(OR4_389_Y), .C(OR4_85_Y), .D(
        OR4_1329_Y), .Y(OR4_699_Y));
    OR4 OR4_12 (.A(\SB_CORRECT[0] ), .B(\SB_CORRECT[1] ), .C(
        \SB_CORRECT[2] ), .D(\SB_CORRECT[3] ), .Y(OR4_12_Y));
    OR4 OR4_978 (.A(OR4_431_Y), .B(OR4_911_Y), .C(OR4_1375_Y), .D(
        OR4_365_Y), .Y(OR4_978_Y));
    CFG3 #( .INIT(8'h2) )  CFG3_12 (.A(W_EN), .B(W_ADDR[15]), .C(
        W_ADDR[14]), .Y(CFG3_12_Y));
    AND4 \AND4SB_CORRECT[105]  (.A(sel_SB_CORRECT_NG[105] ), .B(
        \BLKY2_pipe[26] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[105] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%31%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R31C0 (.A_DOUT({
        nc888, nc889, nc890, nc891, nc892,int_R_DATA_TEMPR31[31] , 
       int_R_DATA_TEMPR31[30] ,int_R_DATA_TEMPR31[29] , 
       int_R_DATA_TEMPR31[28] ,int_R_DATA_TEMPR31[27] , 
       int_R_DATA_TEMPR31[26] ,int_R_DATA_TEMPR31[25] , 
       int_R_DATA_TEMPR31[24] ,int_R_DATA_TEMPR31[23] , 
       int_R_DATA_TEMPR31[22] ,int_R_DATA_TEMPR31[21] , 
       int_R_DATA_TEMPR31[20] ,int_R_DATA_TEMPR31[19] , 
       int_R_DATA_TEMPR31[18] ,int_R_DATA_TEMPR31[17] }), .B_DOUT({nc893, 
        nc894, nc895,int_R_DATA_TEMPR31[16] ,int_R_DATA_TEMPR31[15] , 
       int_R_DATA_TEMPR31[14] ,int_R_DATA_TEMPR31[13] , 
       int_R_DATA_TEMPR31[12] ,int_R_DATA_TEMPR31[11] , 
       int_R_DATA_TEMPR31[10] ,int_R_DATA_TEMPR31[9] ,int_R_DATA_TEMPR31[8] , 
       int_R_DATA_TEMPR31[7] ,int_R_DATA_TEMPR31[6] ,int_R_DATA_TEMPR31[5] , 
       int_R_DATA_TEMPR31[4] ,int_R_DATA_TEMPR31[3] ,int_R_DATA_TEMPR31[2] , 
       int_R_DATA_TEMPR31[1] ,int_R_DATA_TEMPR31[0] }), .DB_DETECT( int_DB_DETECT_NG[31] ), .SB_CORRECT(int_SB_CORRECT_NG[31] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[31] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[7] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[7] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_583 (.A(sel_R_DATA_TEMPR0[31] ), .B(sel_R_DATA_TEMPR1[31] ), .C(sel_R_DATA_TEMPR2[31] ), .D(sel_R_DATA_TEMPR3[31] ), .Y(OR4_583_Y));
    OR4 OR4_412 (.A(sel_R_DATA_TEMPR68[21] ), .B(sel_R_DATA_TEMPR69[21] ), 
        .C(sel_R_DATA_TEMPR70[21] ), .D(sel_R_DATA_TEMPR71[21] ), .Y(
        OR4_412_Y));
    OR4 OR4_1035 (.A(sel_R_DATA_TEMPR40[25] ), .B(sel_R_DATA_TEMPR41[25] ), 
        .C(sel_R_DATA_TEMPR42[25] ), .D(sel_R_DATA_TEMPR43[25] ), .Y(
        OR4_1035_Y));
    AND4 \AND4SB_CORRECT[44]  (.A(sel_SB_CORRECT_NG[44] ), .B(
        \BLKY2_pipe[11] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[44] ));
    OR4 OR4_296 (.A(\SB_CORRECT[124] ), .B(\SB_CORRECT[125] ), 
        .C(\SB_CORRECT[126] ), .D(\SB_CORRECT[127] ), .Y(
        OR4_296_Y));
    AND4 \AND4SB_CORRECT[114]  (.A(sel_SB_CORRECT_NG[114] ), .B(
        \BLKY2_pipe[28] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[114] ));
    OR4 OR4_1121 (.A(sel_R_DATA_TEMPR120[31] ), .B(sel_R_DATA_TEMPR121[31] ), 
        .C(sel_R_DATA_TEMPR122[31] ), .D(sel_R_DATA_TEMPR123[31] ), .Y(
        OR4_1121_Y));
    OR4 OR4_1056 (.A(sel_R_DATA_TEMPR96[2] ), .B(sel_R_DATA_TEMPR97[2] ), .C(sel_R_DATA_TEMPR98[2] ), .D(sel_R_DATA_TEMPR99[2] ), .Y(OR4_1056_Y));
    OR4 OR4_419 (.A(sel_R_DATA_TEMPR100[11] ), .B(sel_R_DATA_TEMPR101[11] ), 
        .C(sel_R_DATA_TEMPR102[11] ), .D(sel_R_DATA_TEMPR103[11] ), .Y(
        OR4_419_Y));
    OR4 OR4_251 (.A(sel_R_DATA_TEMPR56[15] ), .B(sel_R_DATA_TEMPR57[15] ), 
        .C(sel_R_DATA_TEMPR58[15] ), .D(sel_R_DATA_TEMPR59[15] ), .Y(
        OR4_251_Y));
    OR4 OR4_79 (.A(sel_R_DATA_TEMPR112[14] ), .B(sel_R_DATA_TEMPR113[14] ), 
        .C(sel_R_DATA_TEMPR114[14] ), .D(sel_R_DATA_TEMPR115[14] ), .Y(
        OR4_79_Y));
    AND4 \AND4DB_DETECT[90]  (.A(sel_DB_DETECT_NG[90] ), .B(
        \BLKY2_pipe[22] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[90] ));
    CFG3 #( .INIT(8'h40) )  CFG3_19 (.A(R_ADDR[13]), .B(R_ADDR[12]), 
        .C(R_ADDR[11]), .Y(CFG3_19_Y));
    OR4 OR4_139 (.A(sel_R_DATA_TEMPR48[23] ), .B(sel_R_DATA_TEMPR49[23] ), 
        .C(sel_R_DATA_TEMPR50[23] ), .D(sel_R_DATA_TEMPR51[23] ), .Y(
        OR4_139_Y));
    AND4 \AND4SB_CORRECT[9]  (.A(sel_SB_CORRECT_NG[9] ), .B(
        \BLKY2_pipe[2] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \SB_CORRECT[9] ));
    OR4 OR4_116 (.A(sel_R_DATA_TEMPR108[8] ), .B(sel_R_DATA_TEMPR109[8] ), 
        .C(sel_R_DATA_TEMPR110[8] ), .D(sel_R_DATA_TEMPR111[8] ), .Y(
        OR4_116_Y));
    OR4 OR4_1182 (.A(sel_R_DATA_TEMPR48[0] ), .B(sel_R_DATA_TEMPR49[0] ), .C(sel_R_DATA_TEMPR50[0] ), .D(sel_R_DATA_TEMPR51[0] ), .Y(OR4_1182_Y));
    OR4 OR4_608 (.A(sel_R_DATA_TEMPR104[20] ), .B(sel_R_DATA_TEMPR105[20] ), 
        .C(sel_R_DATA_TEMPR106[20] ), .D(sel_R_DATA_TEMPR107[20] ), .Y(
        OR4_608_Y));
    OR4 OR4_144 (.A(sel_R_DATA_TEMPR72[19] ), .B(sel_R_DATA_TEMPR73[19] ), 
        .C(sel_R_DATA_TEMPR74[19] ), .D(sel_R_DATA_TEMPR75[19] ), .Y(
        OR4_144_Y));
    AND4 \AND4DB_DETECT[5]  (.A(sel_DB_DETECT_NG[5] ), .B(
        \BLKY2_pipe[1] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[5] ));
    OR4 OR4_694 (.A(sel_R_DATA_TEMPR56[3] ), .B(sel_R_DATA_TEMPR57[3] ), .C(sel_R_DATA_TEMPR58[3] ), .D(sel_R_DATA_TEMPR59[3] ), .Y(OR4_694_Y));
    OR4 OR4_1351 (.A(OR4_1004_Y), .B(OR4_1243_Y), .C(OR4_797_Y), .D(
        OR4_576_Y), .Y(OR4_1351_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%101%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R101C0 (.A_DOUT({
        nc896, nc897, nc898, nc899, nc900,int_R_DATA_TEMPR101[31] , 
       int_R_DATA_TEMPR101[30] ,int_R_DATA_TEMPR101[29] , 
       int_R_DATA_TEMPR101[28] ,int_R_DATA_TEMPR101[27] , 
       int_R_DATA_TEMPR101[26] ,int_R_DATA_TEMPR101[25] , 
       int_R_DATA_TEMPR101[24] ,int_R_DATA_TEMPR101[23] , 
       int_R_DATA_TEMPR101[22] ,int_R_DATA_TEMPR101[21] , 
       int_R_DATA_TEMPR101[20] ,int_R_DATA_TEMPR101[19] , 
       int_R_DATA_TEMPR101[18] ,int_R_DATA_TEMPR101[17] }), .B_DOUT({nc901, 
        nc902, nc903,int_R_DATA_TEMPR101[16] ,int_R_DATA_TEMPR101[15] , 
       int_R_DATA_TEMPR101[14] ,int_R_DATA_TEMPR101[13] , 
       int_R_DATA_TEMPR101[12] ,int_R_DATA_TEMPR101[11] , 
       int_R_DATA_TEMPR101[10] ,int_R_DATA_TEMPR101[9] , 
       int_R_DATA_TEMPR101[8] ,int_R_DATA_TEMPR101[7] , 
       int_R_DATA_TEMPR101[6] ,int_R_DATA_TEMPR101[5] , 
       int_R_DATA_TEMPR101[4] ,int_R_DATA_TEMPR101[3] , 
       int_R_DATA_TEMPR101[2] ,int_R_DATA_TEMPR101[1] , 
       int_R_DATA_TEMPR101[0] }), .DB_DETECT(int_DB_DETECT_NG[101] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[101] ), .ACCESS_BUSY(
        ACCESS_BUSY[101] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[25] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[25] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4DB_DETECT[60]  (.A(sel_DB_DETECT_NG[60] ), .B(
        \BLKY2_pipe[15] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[60] ));
    OR4 OR4_678 (.A(\DB_DETECT[108] ), .B(\DB_DETECT[109] ), .C(
        \DB_DETECT[110] ), .D(\DB_DETECT[111] ), .Y(OR4_678_Y));
    OR4 OR4_602 (.A(OR4_593_Y), .B(OR4_382_Y), .C(OR4_130_Y), .D(
        OR4_393_Y), .Y(OR4_602_Y));
    OR4 OR4_552 (.A(OR4_343_Y), .B(OR4_979_Y), .C(OR4_60_Y), .D(
        OR4_926_Y), .Y(OR4_552_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[25]  (.A(CFG3_8_Y), .B(CFG3_7_Y)
        , .Y(\BLKX2[25] ));
    AND4 \AND4SB_CORRECT[6]  (.A(sel_SB_CORRECT_NG[6] ), .B(
        \BLKY2_pipe[1] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[6] ));
    OR4 OR4_931 (.A(sel_R_DATA_TEMPR36[13] ), .B(sel_R_DATA_TEMPR37[13] ), 
        .C(sel_R_DATA_TEMPR38[13] ), .D(sel_R_DATA_TEMPR39[13] ), .Y(
        OR4_931_Y));
    OR4 OR4_943 (.A(sel_R_DATA_TEMPR4[20] ), .B(sel_R_DATA_TEMPR5[20] ), .C(sel_R_DATA_TEMPR6[20] ), .D(sel_R_DATA_TEMPR7[20] ), .Y(OR4_943_Y));
    OR4 OR4_220 (.A(sel_R_DATA_TEMPR32[26] ), .B(sel_R_DATA_TEMPR33[26] ), 
        .C(sel_R_DATA_TEMPR34[26] ), .D(sel_R_DATA_TEMPR35[26] ), .Y(
        OR4_220_Y));
    OR4 OR4_1273 (.A(sel_R_DATA_TEMPR60[4] ), .B(sel_R_DATA_TEMPR61[4] ), .C(sel_R_DATA_TEMPR62[4] ), .D(sel_R_DATA_TEMPR63[4] ), .Y(OR4_1273_Y));
    AND4 \AND4DB_DETECT[89]  (.A(sel_DB_DETECT_NG[89] ), .B(
        \BLKY2_pipe[22] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[89] ));
    OR4 OR4_672 (.A(sel_R_DATA_TEMPR8[31] ), .B(sel_R_DATA_TEMPR9[31] ), .C(sel_R_DATA_TEMPR10[31] ), .D(sel_R_DATA_TEMPR11[31] ), .Y(OR4_672_Y));
    OR4 OR4_527 (.A(sel_R_DATA_TEMPR40[6] ), .B(sel_R_DATA_TEMPR41[6] ), .C(sel_R_DATA_TEMPR42[6] ), .D(sel_R_DATA_TEMPR43[6] ), .Y(OR4_527_Y));
    OR4 OR4_318 (.A(sel_R_DATA_TEMPR104[5] ), .B(sel_R_DATA_TEMPR105[5] ), 
        .C(sel_R_DATA_TEMPR106[5] ), .D(sel_R_DATA_TEMPR107[5] ), .Y(
        OR4_318_Y));
    OR2 OR2_10 (.A(\DB_DETECT[84] ), .B(\DB_DETECT[85] ), .Y(
        OR2_10_Y));
    AND4 \AND4DB_DETECT[16]  (.A(sel_DB_DETECT_NG[16] ), .B(
        \BLKY2_pipe[4] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[16] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%117%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R117C0 (.A_DOUT({
        nc904, nc905, nc906, nc907, nc908,int_R_DATA_TEMPR117[31] , 
       int_R_DATA_TEMPR117[30] ,int_R_DATA_TEMPR117[29] , 
       int_R_DATA_TEMPR117[28] ,int_R_DATA_TEMPR117[27] , 
       int_R_DATA_TEMPR117[26] ,int_R_DATA_TEMPR117[25] , 
       int_R_DATA_TEMPR117[24] ,int_R_DATA_TEMPR117[23] , 
       int_R_DATA_TEMPR117[22] ,int_R_DATA_TEMPR117[21] , 
       int_R_DATA_TEMPR117[20] ,int_R_DATA_TEMPR117[19] , 
       int_R_DATA_TEMPR117[18] ,int_R_DATA_TEMPR117[17] }), .B_DOUT({nc909, 
        nc910, nc911,int_R_DATA_TEMPR117[16] ,int_R_DATA_TEMPR117[15] , 
       int_R_DATA_TEMPR117[14] ,int_R_DATA_TEMPR117[13] , 
       int_R_DATA_TEMPR117[12] ,int_R_DATA_TEMPR117[11] , 
       int_R_DATA_TEMPR117[10] ,int_R_DATA_TEMPR117[9] , 
       int_R_DATA_TEMPR117[8] ,int_R_DATA_TEMPR117[7] , 
       int_R_DATA_TEMPR117[6] ,int_R_DATA_TEMPR117[5] , 
       int_R_DATA_TEMPR117[4] ,int_R_DATA_TEMPR117[3] , 
       int_R_DATA_TEMPR117[2] ,int_R_DATA_TEMPR117[1] , 
       int_R_DATA_TEMPR117[0] }), .DB_DETECT(int_DB_DETECT_NG[117] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[117] ), .ACCESS_BUSY(
        ACCESS_BUSY[117] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[29] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), .A_DIN({GND, 
        GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[29] , \BLKX1[0] , W_ADDR[9]}), .B_CLK(
        CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_846 (.A(OR4_1195_Y), .B(OR4_66_Y), .C(OR4_970_Y), .D(
        OR4_317_Y), .Y(OR4_846_Y));
    OR4 OR4_741 (.A(sel_R_DATA_TEMPR4[7] ), .B(sel_R_DATA_TEMPR5[7] ), .C(sel_R_DATA_TEMPR6[7] ), .D(sel_R_DATA_TEMPR7[7] ), .Y(OR4_741_Y));
    AND4 \AND4DB_DETECT[11]  (.A(sel_DB_DETECT_NG[11] ), .B(
        \BLKY2_pipe[2] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[11] ));
    OR4 OR4_1012 (.A(sel_R_DATA_TEMPR8[3] ), .B(sel_R_DATA_TEMPR9[3] ), .C(sel_R_DATA_TEMPR10[3] ), .D(sel_R_DATA_TEMPR11[3] ), .Y(OR4_1012_Y));
    OR4 \OR4_R_DATA[3]  (.A(OR4_331_Y), .B(OR4_710_Y), .C(OR4_599_Y), 
        .D(OR4_706_Y), .Y(R_DATA[3]));
    AND4 \AND4DB_DETECT[105]  (.A(sel_DB_DETECT_NG[105] ), .B(
        \BLKY2_pipe[26] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[105] ));
    OR2 OR2_17 (.A(sel_R_DATA_TEMPR84[9] ), .B(sel_R_DATA_TEMPR85[9] ), .Y(
        OR2_17_Y));
    OR4 OR4_666 (.A(sel_R_DATA_TEMPR120[9] ), .B(sel_R_DATA_TEMPR121[9] ), 
        .C(sel_R_DATA_TEMPR122[9] ), .D(sel_R_DATA_TEMPR123[9] ), .Y(
        OR4_666_Y));
    OR4 OR4_629 (.A(sel_R_DATA_TEMPR80[10] ), .B(sel_R_DATA_TEMPR81[10] ), 
        .C(sel_R_DATA_TEMPR82[10] ), .D(sel_R_DATA_TEMPR83[10] ), .Y(
        OR4_629_Y));
    OR4 OR4_1025 (.A(sel_R_DATA_TEMPR64[1] ), .B(sel_R_DATA_TEMPR65[1] ), .C(sel_R_DATA_TEMPR66[1] ), .D(sel_R_DATA_TEMPR67[1] ), .Y(OR4_1025_Y));
    OR4 OR4_554 (.A(sel_R_DATA_TEMPR116[5] ), .B(sel_R_DATA_TEMPR117[5] ), 
        .C(sel_R_DATA_TEMPR118[5] ), .D(sel_R_DATA_TEMPR119[5] ), .Y(
        OR4_554_Y));
    AND4 \AND4SB_CORRECT[71]  (.A(sel_SB_CORRECT_NG[71] ), .B(
        \BLKY2_pipe[17] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[71] ));
    OR4 OR4_952 (.A(sel_R_DATA_TEMPR92[15] ), .B(sel_R_DATA_TEMPR93[15] ), 
        .C(sel_R_DATA_TEMPR94[15] ), .D(sel_R_DATA_TEMPR95[15] ), .Y(
        OR4_952_Y));
    OR4 OR4_546 (.A(sel_R_DATA_TEMPR120[19] ), .B(sel_R_DATA_TEMPR121[19] ), 
        .C(sel_R_DATA_TEMPR122[19] ), .D(sel_R_DATA_TEMPR123[19] ), .Y(
        OR4_546_Y));
    OR4 OR4_226 (.A(sel_R_DATA_TEMPR0[18] ), .B(sel_R_DATA_TEMPR1[18] ), .C(sel_R_DATA_TEMPR2[18] ), .D(sel_R_DATA_TEMPR3[18] ), .Y(OR4_226_Y));
    OR4 OR4_119 (.A(sel_R_DATA_TEMPR112[23] ), .B(sel_R_DATA_TEMPR113[23] ), 
        .C(sel_R_DATA_TEMPR114[23] ), .D(sel_R_DATA_TEMPR115[23] ), .Y(
        OR4_119_Y));
    AND4 \AND4DB_DETECT[124]  (.A(sel_DB_DETECT_NG[124] ), .B(
        \BLKY2_pipe[31] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[124] ));
    OR4 OR4_1047 (.A(OR4_1364_Y), .B(OR4_184_Y), .C(OR4_1157_Y), .D(
        OR4_927_Y), .Y(OR4_1047_Y));
    OR4 OR4_805 (.A(sel_R_DATA_TEMPR44[27] ), .B(sel_R_DATA_TEMPR45[27] ), 
        .C(sel_R_DATA_TEMPR46[27] ), .D(sel_R_DATA_TEMPR47[27] ), .Y(
        OR4_805_Y));
    OR4 OR4_1179 (.A(sel_R_DATA_TEMPR112[4] ), .B(sel_R_DATA_TEMPR113[4] ), 
        .C(sel_R_DATA_TEMPR114[4] ), .D(sel_R_DATA_TEMPR115[4] ), .Y(
        OR4_1179_Y));
    OR4 OR4_72 (.A(sel_R_DATA_TEMPR116[1] ), .B(sel_R_DATA_TEMPR117[1] ), .C(sel_R_DATA_TEMPR118[1] ), .D(sel_R_DATA_TEMPR119[1] ), .Y(OR4_72_Y));
    AND4 \AND4DB_DETECT[45]  (.A(sel_DB_DETECT_NG[45] ), .B(
        \BLKY2_pipe[11] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[45] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%98%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R98C0 (.A_DOUT({
        nc912, nc913, nc914, nc915, nc916,int_R_DATA_TEMPR98[31] , 
       int_R_DATA_TEMPR98[30] ,int_R_DATA_TEMPR98[29] , 
       int_R_DATA_TEMPR98[28] ,int_R_DATA_TEMPR98[27] , 
       int_R_DATA_TEMPR98[26] ,int_R_DATA_TEMPR98[25] , 
       int_R_DATA_TEMPR98[24] ,int_R_DATA_TEMPR98[23] , 
       int_R_DATA_TEMPR98[22] ,int_R_DATA_TEMPR98[21] , 
       int_R_DATA_TEMPR98[20] ,int_R_DATA_TEMPR98[19] , 
       int_R_DATA_TEMPR98[18] ,int_R_DATA_TEMPR98[17] }), .B_DOUT({nc917, 
        nc918, nc919,int_R_DATA_TEMPR98[16] ,int_R_DATA_TEMPR98[15] , 
       int_R_DATA_TEMPR98[14] ,int_R_DATA_TEMPR98[13] , 
       int_R_DATA_TEMPR98[12] ,int_R_DATA_TEMPR98[11] , 
       int_R_DATA_TEMPR98[10] ,int_R_DATA_TEMPR98[9] ,int_R_DATA_TEMPR98[8] , 
       int_R_DATA_TEMPR98[7] ,int_R_DATA_TEMPR98[6] ,int_R_DATA_TEMPR98[5] , 
       int_R_DATA_TEMPR98[4] ,int_R_DATA_TEMPR98[3] ,int_R_DATA_TEMPR98[2] , 
       int_R_DATA_TEMPR98[1] ,int_R_DATA_TEMPR98[0] }), .DB_DETECT( int_DB_DETECT_NG[98] ), .SB_CORRECT(int_SB_CORRECT_NG[98] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[98] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[24] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[24] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1130 (.A(sel_R_DATA_TEMPR28[30] ), .B(sel_R_DATA_TEMPR29[30] ), 
        .C(sel_R_DATA_TEMPR30[30] ), .D(sel_R_DATA_TEMPR31[30] ), .Y(
        OR4_1130_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%95%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R95C0 (.A_DOUT({
        nc920, nc921, nc922, nc923, nc924,int_R_DATA_TEMPR95[31] , 
       int_R_DATA_TEMPR95[30] ,int_R_DATA_TEMPR95[29] , 
       int_R_DATA_TEMPR95[28] ,int_R_DATA_TEMPR95[27] , 
       int_R_DATA_TEMPR95[26] ,int_R_DATA_TEMPR95[25] , 
       int_R_DATA_TEMPR95[24] ,int_R_DATA_TEMPR95[23] , 
       int_R_DATA_TEMPR95[22] ,int_R_DATA_TEMPR95[21] , 
       int_R_DATA_TEMPR95[20] ,int_R_DATA_TEMPR95[19] , 
       int_R_DATA_TEMPR95[18] ,int_R_DATA_TEMPR95[17] }), .B_DOUT({nc925, 
        nc926, nc927,int_R_DATA_TEMPR95[16] ,int_R_DATA_TEMPR95[15] , 
       int_R_DATA_TEMPR95[14] ,int_R_DATA_TEMPR95[13] , 
       int_R_DATA_TEMPR95[12] ,int_R_DATA_TEMPR95[11] , 
       int_R_DATA_TEMPR95[10] ,int_R_DATA_TEMPR95[9] ,int_R_DATA_TEMPR95[8] , 
       int_R_DATA_TEMPR95[7] ,int_R_DATA_TEMPR95[6] ,int_R_DATA_TEMPR95[5] , 
       int_R_DATA_TEMPR95[4] ,int_R_DATA_TEMPR95[3] ,int_R_DATA_TEMPR95[2] , 
       int_R_DATA_TEMPR95[1] ,int_R_DATA_TEMPR95[0] }), .DB_DETECT( int_DB_DETECT_NG[95] ), .SB_CORRECT(int_SB_CORRECT_NG[95] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[95] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[23] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[23] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_875 (.A(OR4_742_Y), .B(OR4_1000_Y), .C(OR4_536_Y), .D(
        OR4_1273_Y), .Y(OR4_875_Y));
    OR4 OR4_735 (.A(sel_R_DATA_TEMPR76[3] ), .B(sel_R_DATA_TEMPR77[3] ), .C(sel_R_DATA_TEMPR78[3] ), .D(sel_R_DATA_TEMPR79[3] ), .Y(OR4_735_Y));
    OR4 OR4_637 (.A(sel_R_DATA_TEMPR100[29] ), .B(sel_R_DATA_TEMPR101[29] ), 
        .C(sel_R_DATA_TEMPR102[29] ), .D(sel_R_DATA_TEMPR103[29] ), .Y(
        OR4_637_Y));
    AND4 \AND4DB_DETECT[115]  (.A(sel_DB_DETECT_NG[115] ), .B(
        \BLKY2_pipe[28] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[115] ));
    AND4 \AND4DB_DETECT[34]  (.A(sel_DB_DETECT_NG[34] ), .B(
        \BLKY2_pipe[8] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[34] ));
    OR4 OR4_736 (.A(sel_R_DATA_TEMPR20[0] ), .B(sel_R_DATA_TEMPR21[0] ), .C(sel_R_DATA_TEMPR22[0] ), .D(sel_R_DATA_TEMPR23[0] ), .Y(OR4_736_Y));
    OR4 OR4_624 (.A(sel_R_DATA_TEMPR8[13] ), .B(sel_R_DATA_TEMPR9[13] ), .C(sel_R_DATA_TEMPR10[13] ), .D(sel_R_DATA_TEMPR11[13] ), .Y(OR4_624_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[30]  (.A(CFG3_10_Y), .B(
        CFG3_7_Y), .Y(\BLKX2[30] ));
    OR4 OR4_351 (.A(sel_R_DATA_TEMPR60[1] ), .B(sel_R_DATA_TEMPR61[1] ), .C(sel_R_DATA_TEMPR62[1] ), .D(sel_R_DATA_TEMPR63[1] ), .Y(OR4_351_Y));
    OR2 OR2_28 (.A(sel_R_DATA_TEMPR84[17] ), .B(sel_R_DATA_TEMPR85[17] ), .Y(
        OR2_28_Y));
    OR4 OR4_911 (.A(sel_R_DATA_TEMPR36[5] ), .B(sel_R_DATA_TEMPR37[5] ), .C(sel_R_DATA_TEMPR38[5] ), .D(sel_R_DATA_TEMPR39[5] ), .Y(OR4_911_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%63%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R63C0 (.A_DOUT({
        nc928, nc929, nc930, nc931, nc932,int_R_DATA_TEMPR63[31] , 
       int_R_DATA_TEMPR63[30] ,int_R_DATA_TEMPR63[29] , 
       int_R_DATA_TEMPR63[28] ,int_R_DATA_TEMPR63[27] , 
       int_R_DATA_TEMPR63[26] ,int_R_DATA_TEMPR63[25] , 
       int_R_DATA_TEMPR63[24] ,int_R_DATA_TEMPR63[23] , 
       int_R_DATA_TEMPR63[22] ,int_R_DATA_TEMPR63[21] , 
       int_R_DATA_TEMPR63[20] ,int_R_DATA_TEMPR63[19] , 
       int_R_DATA_TEMPR63[18] ,int_R_DATA_TEMPR63[17] }), .B_DOUT({nc933, 
        nc934, nc935,int_R_DATA_TEMPR63[16] ,int_R_DATA_TEMPR63[15] , 
       int_R_DATA_TEMPR63[14] ,int_R_DATA_TEMPR63[13] , 
       int_R_DATA_TEMPR63[12] ,int_R_DATA_TEMPR63[11] , 
       int_R_DATA_TEMPR63[10] ,int_R_DATA_TEMPR63[9] ,int_R_DATA_TEMPR63[8] , 
       int_R_DATA_TEMPR63[7] ,int_R_DATA_TEMPR63[6] ,int_R_DATA_TEMPR63[5] , 
       int_R_DATA_TEMPR63[4] ,int_R_DATA_TEMPR63[3] ,int_R_DATA_TEMPR63[2] , 
       int_R_DATA_TEMPR63[1] ,int_R_DATA_TEMPR63[0] }), .DB_DETECT( int_DB_DETECT_NG[63] ), .SB_CORRECT(int_SB_CORRECT_NG[63] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[63] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[15] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[15] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4SB_CORRECT[10]  (.A(sel_SB_CORRECT_NG[10] ), .B(
        \BLKY2_pipe[2] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[10] ));
    OR4 OR4_1365 (.A(sel_R_DATA_TEMPR16[23] ), .B(sel_R_DATA_TEMPR17[23] ), 
        .C(sel_R_DATA_TEMPR18[23] ), .D(sel_R_DATA_TEMPR19[23] ), .Y(
        OR4_1365_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[9]  (.D(\BLKY2[9] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[9] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%124%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R124C0 (.A_DOUT({
        nc936, nc937, nc938, nc939, nc940,int_R_DATA_TEMPR124[31] , 
       int_R_DATA_TEMPR124[30] ,int_R_DATA_TEMPR124[29] , 
       int_R_DATA_TEMPR124[28] ,int_R_DATA_TEMPR124[27] , 
       int_R_DATA_TEMPR124[26] ,int_R_DATA_TEMPR124[25] , 
       int_R_DATA_TEMPR124[24] ,int_R_DATA_TEMPR124[23] , 
       int_R_DATA_TEMPR124[22] ,int_R_DATA_TEMPR124[21] , 
       int_R_DATA_TEMPR124[20] ,int_R_DATA_TEMPR124[19] , 
       int_R_DATA_TEMPR124[18] ,int_R_DATA_TEMPR124[17] }), .B_DOUT({nc941, 
        nc942, nc943,int_R_DATA_TEMPR124[16] ,int_R_DATA_TEMPR124[15] , 
       int_R_DATA_TEMPR124[14] ,int_R_DATA_TEMPR124[13] , 
       int_R_DATA_TEMPR124[12] ,int_R_DATA_TEMPR124[11] , 
       int_R_DATA_TEMPR124[10] ,int_R_DATA_TEMPR124[9] , 
       int_R_DATA_TEMPR124[8] ,int_R_DATA_TEMPR124[7] , 
       int_R_DATA_TEMPR124[6] ,int_R_DATA_TEMPR124[5] , 
       int_R_DATA_TEMPR124[4] ,int_R_DATA_TEMPR124[3] , 
       int_R_DATA_TEMPR124[2] ,int_R_DATA_TEMPR124[1] , 
       int_R_DATA_TEMPR124[0] }), .DB_DETECT(int_DB_DETECT_NG[124] ), 
        .SB_CORRECT(int_SB_CORRECT_NG[124] ), .ACCESS_BUSY(
        ACCESS_BUSY[124] ), .A_ADDR({R_ADDR[8], R_ADDR[7], 
        R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], R_ADDR[2], 
        R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), .A_BLK_EN({
        \BLKY2[31] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), .A_DIN({
        GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], W_DATA[29], 
        W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], W_DATA[24], 
        W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], W_DATA[19], 
        W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, VCC}), 
        .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(VCC), 
        .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], W_ADDR[4], 
        W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, GND, GND, GND, 
        GND}), .B_BLK_EN({\BLKX2[31] , \BLKX1[0] , \BLKX0[0] }), 
        .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], W_DATA[15], 
        W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], W_DATA[10], 
        W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], W_DATA[5], 
        W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], W_DATA[0]}), 
        .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_450 (.A(sel_R_DATA_TEMPR116[19] ), .B(sel_R_DATA_TEMPR117[19] ), 
        .C(sel_R_DATA_TEMPR118[19] ), .D(sel_R_DATA_TEMPR119[19] ), .Y(
        OR4_450_Y));
    OR4 \OR4_R_DATA[25]  (.A(OR4_1086_Y), .B(OR4_367_Y), .C(OR4_894_Y), 
        .D(OR4_510_Y), .Y(R_DATA[25]));
    OR4 OR4_283 (.A(OR4_747_Y), .B(OR4_594_Y), .C(OR4_99_Y), .D(
        OR4_529_Y), .Y(OR4_283_Y));
    OR4 OR4_96 (.A(sel_R_DATA_TEMPR52[1] ), .B(sel_R_DATA_TEMPR53[1] ), .C(sel_R_DATA_TEMPR54[1] ), .D(sel_R_DATA_TEMPR55[1] ), .Y(OR4_96_Y));
    OR4 OR4_1209 (.A(sel_R_DATA_TEMPR80[14] ), .B(sel_R_DATA_TEMPR81[14] ), 
        .C(sel_R_DATA_TEMPR82[14] ), .D(sel_R_DATA_TEMPR83[14] ), .Y(
        OR4_1209_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%52%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R52C0 (.A_DOUT({
        nc944, nc945, nc946, nc947, nc948,int_R_DATA_TEMPR52[31] , 
       int_R_DATA_TEMPR52[30] ,int_R_DATA_TEMPR52[29] , 
       int_R_DATA_TEMPR52[28] ,int_R_DATA_TEMPR52[27] , 
       int_R_DATA_TEMPR52[26] ,int_R_DATA_TEMPR52[25] , 
       int_R_DATA_TEMPR52[24] ,int_R_DATA_TEMPR52[23] , 
       int_R_DATA_TEMPR52[22] ,int_R_DATA_TEMPR52[21] , 
       int_R_DATA_TEMPR52[20] ,int_R_DATA_TEMPR52[19] , 
       int_R_DATA_TEMPR52[18] ,int_R_DATA_TEMPR52[17] }), .B_DOUT({nc949, 
        nc950, nc951,int_R_DATA_TEMPR52[16] ,int_R_DATA_TEMPR52[15] , 
       int_R_DATA_TEMPR52[14] ,int_R_DATA_TEMPR52[13] , 
       int_R_DATA_TEMPR52[12] ,int_R_DATA_TEMPR52[11] , 
       int_R_DATA_TEMPR52[10] ,int_R_DATA_TEMPR52[9] ,int_R_DATA_TEMPR52[8] , 
       int_R_DATA_TEMPR52[7] ,int_R_DATA_TEMPR52[6] ,int_R_DATA_TEMPR52[5] , 
       int_R_DATA_TEMPR52[4] ,int_R_DATA_TEMPR52[3] ,int_R_DATA_TEMPR52[2] , 
       int_R_DATA_TEMPR52[1] ,int_R_DATA_TEMPR52[0] }), .DB_DETECT( int_DB_DETECT_NG[52] ), .SB_CORRECT(int_SB_CORRECT_NG[52] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[52] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[13] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[13] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    CFG3 #( .INIT(8'h8) )  CFG3_17 (.A(W_EN), .B(W_ADDR[15]), .C(
        W_ADDR[14]), .Y(CFG3_17_Y));
    OR4 OR4_1330 (.A(sel_R_DATA_TEMPR124[1] ), .B(sel_R_DATA_TEMPR125[1] ), 
        .C(sel_R_DATA_TEMPR126[1] ), .D(sel_R_DATA_TEMPR127[1] ), .Y(
        OR4_1330_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%87%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R87C0 (.A_DOUT({
        nc952, nc953, nc954, nc955, nc956,int_R_DATA_TEMPR87[31] , 
       int_R_DATA_TEMPR87[30] ,int_R_DATA_TEMPR87[29] , 
       int_R_DATA_TEMPR87[28] ,int_R_DATA_TEMPR87[27] , 
       int_R_DATA_TEMPR87[26] ,int_R_DATA_TEMPR87[25] , 
       int_R_DATA_TEMPR87[24] ,int_R_DATA_TEMPR87[23] , 
       int_R_DATA_TEMPR87[22] ,int_R_DATA_TEMPR87[21] , 
       int_R_DATA_TEMPR87[20] ,int_R_DATA_TEMPR87[19] , 
       int_R_DATA_TEMPR87[18] ,int_R_DATA_TEMPR87[17] }), .B_DOUT({nc957, 
        nc958, nc959,int_R_DATA_TEMPR87[16] ,int_R_DATA_TEMPR87[15] , 
       int_R_DATA_TEMPR87[14] ,int_R_DATA_TEMPR87[13] , 
       int_R_DATA_TEMPR87[12] ,int_R_DATA_TEMPR87[11] , 
       int_R_DATA_TEMPR87[10] ,int_R_DATA_TEMPR87[9] ,int_R_DATA_TEMPR87[8] , 
       int_R_DATA_TEMPR87[7] ,int_R_DATA_TEMPR87[6] ,int_R_DATA_TEMPR87[5] , 
       int_R_DATA_TEMPR87[4] ,int_R_DATA_TEMPR87[3] ,int_R_DATA_TEMPR87[2] , 
       int_R_DATA_TEMPR87[1] ,int_R_DATA_TEMPR87[0] }), .DB_DETECT( int_DB_DETECT_NG[87] ), .SB_CORRECT(int_SB_CORRECT_NG[87] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[87] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[21] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[21] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1176 (.A(sel_R_DATA_TEMPR32[22] ), .B(sel_R_DATA_TEMPR33[22] ), 
        .C(sel_R_DATA_TEMPR34[22] ), .D(sel_R_DATA_TEMPR35[22] ), .Y(
        OR4_1176_Y));
    OR4 OR4_548 (.A(sel_R_DATA_TEMPR108[23] ), .B(sel_R_DATA_TEMPR109[23] ), 
        .C(sel_R_DATA_TEMPR110[23] ), .D(sel_R_DATA_TEMPR111[23] ), .Y(
        OR4_548_Y));
    OR4 OR4_1152 (.A(sel_R_DATA_TEMPR20[20] ), .B(sel_R_DATA_TEMPR21[20] ), 
        .C(sel_R_DATA_TEMPR22[20] ), .D(sel_R_DATA_TEMPR23[20] ), .Y(
        OR4_1152_Y));
    OR4 OR4_54 (.A(OR4_442_Y), .B(OR4_302_Y), .C(OR4_403_Y), .D(
        OR4_80_Y), .Y(OR4_54_Y));
    AND4 \AND4DB_DETECT[73]  (.A(sel_DB_DETECT_NG[73] ), .B(
        \BLKY2_pipe[18] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[73] ));
    OR4 OR4_988 (.A(OR4_605_Y), .B(OR4_1280_Y), .C(OR4_292_Y), .D(
        OR4_545_Y), .Y(OR4_988_Y));
    OR4 OR4_1271 (.A(sel_R_DATA_TEMPR44[14] ), .B(sel_R_DATA_TEMPR45[14] ), 
        .C(sel_R_DATA_TEMPR46[14] ), .D(sel_R_DATA_TEMPR47[14] ), .Y(
        OR4_1271_Y));
    OR4 OR4_3 (.A(sel_R_DATA_TEMPR116[4] ), .B(sel_R_DATA_TEMPR117[4] ), .C(sel_R_DATA_TEMPR118[4] ), .D(sel_R_DATA_TEMPR119[4] ), .Y(OR4_3_Y));
    AND4 \AND4SB_CORRECT[51]  (.A(sel_SB_CORRECT_NG[51] ), .B(
        \BLKY2_pipe[12] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[51] ));
    DFN1E1 \DFN1E1BLKY2_pipe[14]  (.D(\BLKY2[14] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[14] ));
    OR4 OR4_1178 (.A(sel_R_DATA_TEMPR64[28] ), .B(sel_R_DATA_TEMPR65[28] ), 
        .C(sel_R_DATA_TEMPR66[28] ), .D(sel_R_DATA_TEMPR67[28] ), .Y(
        OR4_1178_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%71%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R71C0 (.A_DOUT({
        nc960, nc961, nc962, nc963, nc964,int_R_DATA_TEMPR71[31] , 
       int_R_DATA_TEMPR71[30] ,int_R_DATA_TEMPR71[29] , 
       int_R_DATA_TEMPR71[28] ,int_R_DATA_TEMPR71[27] , 
       int_R_DATA_TEMPR71[26] ,int_R_DATA_TEMPR71[25] , 
       int_R_DATA_TEMPR71[24] ,int_R_DATA_TEMPR71[23] , 
       int_R_DATA_TEMPR71[22] ,int_R_DATA_TEMPR71[21] , 
       int_R_DATA_TEMPR71[20] ,int_R_DATA_TEMPR71[19] , 
       int_R_DATA_TEMPR71[18] ,int_R_DATA_TEMPR71[17] }), .B_DOUT({nc965, 
        nc966, nc967,int_R_DATA_TEMPR71[16] ,int_R_DATA_TEMPR71[15] , 
       int_R_DATA_TEMPR71[14] ,int_R_DATA_TEMPR71[13] , 
       int_R_DATA_TEMPR71[12] ,int_R_DATA_TEMPR71[11] , 
       int_R_DATA_TEMPR71[10] ,int_R_DATA_TEMPR71[9] ,int_R_DATA_TEMPR71[8] , 
       int_R_DATA_TEMPR71[7] ,int_R_DATA_TEMPR71[6] ,int_R_DATA_TEMPR71[5] , 
       int_R_DATA_TEMPR71[4] ,int_R_DATA_TEMPR71[3] ,int_R_DATA_TEMPR71[2] , 
       int_R_DATA_TEMPR71[1] ,int_R_DATA_TEMPR71[0] }), .DB_DETECT( int_DB_DETECT_NG[71] ), .SB_CORRECT(int_SB_CORRECT_NG[71] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[71] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[17] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[17] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_364 (.A(OR4_949_Y), .B(OR4_234_Y), .C(OR4_623_Y), .D(
        OR4_883_Y), .Y(OR4_364_Y));
    AND4 \AND4DB_DETECT[26]  (.A(sel_DB_DETECT_NG[26] ), .B(
        \BLKY2_pipe[6] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[26] ));
    OR4 OR4_1120 (.A(OR4_1138_Y), .B(OR4_245_Y), .C(OR4_907_Y), .D(
        OR4_1127_Y), .Y(OR4_1120_Y));
    OR4 OR4_606 (.A(OR4_932_Y), .B(OR4_1152_Y), .C(OR4_727_Y), .D(
        OR4_511_Y), .Y(OR4_606_Y));
    AND4 \AND4DB_DETECT[21]  (.A(sel_DB_DETECT_NG[21] ), .B(
        \BLKY2_pipe[5] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[21] ));
    OR4 OR4_715 (.A(sel_R_DATA_TEMPR0[30] ), .B(sel_R_DATA_TEMPR1[30] ), .C(sel_R_DATA_TEMPR2[30] ), .D(sel_R_DATA_TEMPR3[30] ), .Y(OR4_715_Y));
    OR4 OR4_617 (.A(sel_R_DATA_TEMPR96[6] ), .B(sel_R_DATA_TEMPR97[6] ), .C(sel_R_DATA_TEMPR98[6] ), .D(sel_R_DATA_TEMPR99[6] ), .Y(OR4_617_Y));
    OR4 OR4_446 (.A(sel_R_DATA_TEMPR44[2] ), .B(sel_R_DATA_TEMPR45[2] ), .C(sel_R_DATA_TEMPR46[2] ), .D(sel_R_DATA_TEMPR47[2] ), .Y(OR4_446_Y));
    OR4 OR4_161 (.A(sel_R_DATA_TEMPR52[21] ), .B(sel_R_DATA_TEMPR53[21] ), 
        .C(sel_R_DATA_TEMPR54[21] ), .D(sel_R_DATA_TEMPR55[21] ), .Y(
        OR4_161_Y));
    OR4 OR4_716 (.A(sel_R_DATA_TEMPR124[2] ), .B(sel_R_DATA_TEMPR125[2] ), 
        .C(sel_R_DATA_TEMPR126[2] ), .D(sel_R_DATA_TEMPR127[2] ), .Y(
        OR4_716_Y));
    OR4 OR4_676 (.A(sel_R_DATA_TEMPR12[23] ), .B(sel_R_DATA_TEMPR13[23] ), 
        .C(sel_R_DATA_TEMPR14[23] ), .D(sel_R_DATA_TEMPR15[23] ), .Y(
        OR4_676_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[17]  (.D(\BLKY2[17] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[17] ));
    OR4 OR4_1289 (.A(sel_R_DATA_TEMPR40[9] ), .B(sel_R_DATA_TEMPR41[9] ), .C(sel_R_DATA_TEMPR42[9] ), .D(sel_R_DATA_TEMPR43[9] ), .Y(OR4_1289_Y));
    AND4 \AND4DB_DETECT[32]  (.A(sel_DB_DETECT_NG[32] ), .B(
        \BLKY2_pipe[8] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), .Y(
        \DB_DETECT[32] ));
    AND4 \AND4DB_DETECT[98]  (.A(sel_DB_DETECT_NG[98] ), .B(
        \BLKY2_pipe[24] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[98] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[6]  (.A(CFG3_1_Y), .B(CFG3_2_Y), 
        .Y(\BLKY2[6] ));
    OR4 OR4_237 (.A(sel_R_DATA_TEMPR60[9] ), .B(sel_R_DATA_TEMPR61[9] ), .C(sel_R_DATA_TEMPR62[9] ), .D(sel_R_DATA_TEMPR63[9] ), .Y(OR4_237_Y));
    OR4 OR4_898 (.A(OR4_1181_Y), .B(OR4_171_Y), .C(OR4_981_Y), .D(
        OR4_1261_Y), .Y(OR4_898_Y));
    OR4 OR4_688 (.A(sel_R_DATA_TEMPR124[28] ), .B(sel_R_DATA_TEMPR125[28] ), 
        .C(sel_R_DATA_TEMPR126[28] ), .D(sel_R_DATA_TEMPR127[28] ), .Y(
        OR4_688_Y));
    OR4 OR4_137 (.A(sel_R_DATA_TEMPR108[29] ), .B(sel_R_DATA_TEMPR109[29] ), 
        .C(sel_R_DATA_TEMPR110[29] ), .D(sel_R_DATA_TEMPR111[29] ), .Y(
        OR4_137_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%6%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R6C0 (.A_DOUT({
        nc968, nc969, nc970, nc971, nc972,int_R_DATA_TEMPR6[31] , 
       int_R_DATA_TEMPR6[30] ,int_R_DATA_TEMPR6[29] ,int_R_DATA_TEMPR6[28] , 
       int_R_DATA_TEMPR6[27] ,int_R_DATA_TEMPR6[26] ,int_R_DATA_TEMPR6[25] , 
       int_R_DATA_TEMPR6[24] ,int_R_DATA_TEMPR6[23] ,int_R_DATA_TEMPR6[22] , 
       int_R_DATA_TEMPR6[21] ,int_R_DATA_TEMPR6[20] ,int_R_DATA_TEMPR6[19] , 
       int_R_DATA_TEMPR6[18] ,int_R_DATA_TEMPR6[17] }), .B_DOUT({nc973, 
        nc974, nc975,int_R_DATA_TEMPR6[16] ,int_R_DATA_TEMPR6[15] , 
       int_R_DATA_TEMPR6[14] ,int_R_DATA_TEMPR6[13] ,int_R_DATA_TEMPR6[12] , 
       int_R_DATA_TEMPR6[11] ,int_R_DATA_TEMPR6[10] ,int_R_DATA_TEMPR6[9] , 
       int_R_DATA_TEMPR6[8] ,int_R_DATA_TEMPR6[7] ,int_R_DATA_TEMPR6[6] , 
       int_R_DATA_TEMPR6[5] ,int_R_DATA_TEMPR6[4] ,int_R_DATA_TEMPR6[3] , 
       int_R_DATA_TEMPR6[2] ,int_R_DATA_TEMPR6[1] ,int_R_DATA_TEMPR6[0] }), 
        .DB_DETECT(int_DB_DETECT_NG[6] ), .SB_CORRECT( int_SB_CORRECT_NG[6] ), .ACCESS_BUSY(\ACCESS_BUSY[6] ), 
        .A_ADDR({R_ADDR[8], R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], 
        R_ADDR[3], R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, 
        GND}), .A_BLK_EN({\BLKY2[1] , R_ADDR[10], \BLKY0[0] }), .A_CLK(
        CLK), .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[1] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4DB_DETECT[68]  (.A(sel_DB_DETECT_NG[68] ), .B(
        \BLKY2_pipe[17] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[68] ));
    AND4 \AND4SB_CORRECT[7]  (.A(sel_SB_CORRECT_NG[7] ), .B(
        \BLKY2_pipe[1] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), .Y(
        \SB_CORRECT[7] ));
    AND4 \AND4SB_CORRECT[92]  (.A(sel_SB_CORRECT_NG[92] ), .B(
        \BLKY2_pipe[23] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[92] ));
    OR4 OR4_1235 (.A(OR4_404_Y), .B(OR4_661_Y), .C(OR4_858_Y), .D(
        OR4_702_Y), .Y(OR4_1235_Y));
    OR4 OR4_682 (.A(OR4_1284_Y), .B(OR4_157_Y), .C(OR4_361_Y), .D(
        OR4_200_Y), .Y(OR4_682_Y));
    OR4 OR4_342 (.A(OR4_101_Y), .B(OR4_1354_Y), .C(OR4_73_Y), .D(
        OR4_28_Y), .Y(OR4_342_Y));
    OR4 OR4_461 (.A(sel_R_DATA_TEMPR116[21] ), .B(sel_R_DATA_TEMPR117[21] ), 
        .C(sel_R_DATA_TEMPR118[21] ), .D(sel_R_DATA_TEMPR119[21] ), .Y(
        OR4_461_Y));
    OR4 OR4_359 (.A(OR4_1204_Y), .B(OR2_5_Y), .C(sel_R_DATA_TEMPR86[3] ), 
        .D(sel_R_DATA_TEMPR87[3] ), .Y(OR4_359_Y));
    DFN1E1 \DFN1E1BLKY2_pipe[21]  (.D(\BLKY2[21] ), .CLK(CLK), .E(VCC), 
        .Q(\BLKY2_pipe[21] ));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKX2[11]  (.A(CFG3_5_Y), .B(CFG3_4_Y)
        , .Y(\BLKX2[11] ));
    OR4 OR4_14 (.A(sel_R_DATA_TEMPR72[1] ), .B(sel_R_DATA_TEMPR73[1] ), .C(sel_R_DATA_TEMPR74[1] ), .D(sel_R_DATA_TEMPR75[1] ), .Y(OR4_14_Y));
    OR4 OR4_468 (.A(sel_R_DATA_TEMPR20[16] ), .B(sel_R_DATA_TEMPR21[16] ), 
        .C(sel_R_DATA_TEMPR22[16] ), .D(sel_R_DATA_TEMPR23[16] ), .Y(
        OR4_468_Y));
    OR4 OR4_1320 (.A(OR4_888_Y), .B(OR4_598_Y), .C(OR4_376_Y), .D(
        OR4_452_Y), .Y(OR4_1320_Y));
    OR2 OR2_18 (.A(sel_R_DATA_TEMPR84[0] ), .B(sel_R_DATA_TEMPR85[0] ), .Y(
        OR2_18_Y));
    OR4 OR4_1247 (.A(sel_R_DATA_TEMPR112[1] ), .B(sel_R_DATA_TEMPR113[1] ), 
        .C(sel_R_DATA_TEMPR114[1] ), .D(sel_R_DATA_TEMPR115[1] ), .Y(
        OR4_1247_Y));
    OR4 OR4_733 (.A(OR4_1356_Y), .B(OR4_541_Y), .C(OR4_989_Y), .D(
        OR4_1388_Y), .Y(OR4_733_Y));
    OR4 OR4_291 (.A(sel_R_DATA_TEMPR44[9] ), .B(sel_R_DATA_TEMPR45[9] ), .C(sel_R_DATA_TEMPR46[9] ), .D(sel_R_DATA_TEMPR47[9] ), .Y(OR4_291_Y));
    OR4 OR4_234 (.A(sel_R_DATA_TEMPR4[15] ), .B(sel_R_DATA_TEMPR5[15] ), .C(sel_R_DATA_TEMPR6[15] ), .D(sel_R_DATA_TEMPR7[15] ), .Y(OR4_234_Y));
    OR4 OR4_1062 (.A(sel_R_DATA_TEMPR32[17] ), .B(sel_R_DATA_TEMPR33[17] ), 
        .C(sel_R_DATA_TEMPR34[17] ), .D(sel_R_DATA_TEMPR35[17] ), .Y(
        OR4_1062_Y));
    OR4 OR4_90 (.A(\DB_DETECT[120] ), .B(\DB_DETECT[121] ), .C(
        \DB_DETECT[122] ), .D(\DB_DETECT[123] ), .Y(OR4_90_Y));
    OR4 OR4_1344 (.A(sel_R_DATA_TEMPR100[20] ), .B(sel_R_DATA_TEMPR101[20] ), 
        .C(sel_R_DATA_TEMPR102[20] ), .D(sel_R_DATA_TEMPR103[20] ), .Y(
        OR4_1344_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%24%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R24C0 (.A_DOUT({
        nc976, nc977, nc978, nc979, nc980,int_R_DATA_TEMPR24[31] , 
       int_R_DATA_TEMPR24[30] ,int_R_DATA_TEMPR24[29] , 
       int_R_DATA_TEMPR24[28] ,int_R_DATA_TEMPR24[27] , 
       int_R_DATA_TEMPR24[26] ,int_R_DATA_TEMPR24[25] , 
       int_R_DATA_TEMPR24[24] ,int_R_DATA_TEMPR24[23] , 
       int_R_DATA_TEMPR24[22] ,int_R_DATA_TEMPR24[21] , 
       int_R_DATA_TEMPR24[20] ,int_R_DATA_TEMPR24[19] , 
       int_R_DATA_TEMPR24[18] ,int_R_DATA_TEMPR24[17] }), .B_DOUT({nc981, 
        nc982, nc983,int_R_DATA_TEMPR24[16] ,int_R_DATA_TEMPR24[15] , 
       int_R_DATA_TEMPR24[14] ,int_R_DATA_TEMPR24[13] , 
       int_R_DATA_TEMPR24[12] ,int_R_DATA_TEMPR24[11] , 
       int_R_DATA_TEMPR24[10] ,int_R_DATA_TEMPR24[9] ,int_R_DATA_TEMPR24[8] , 
       int_R_DATA_TEMPR24[7] ,int_R_DATA_TEMPR24[6] ,int_R_DATA_TEMPR24[5] , 
       int_R_DATA_TEMPR24[4] ,int_R_DATA_TEMPR24[3] ,int_R_DATA_TEMPR24[2] , 
       int_R_DATA_TEMPR24[1] ,int_R_DATA_TEMPR24[0] }), .DB_DETECT( int_DB_DETECT_NG[24] ), .SB_CORRECT(int_SB_CORRECT_NG[24] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[24] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[6] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[6] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_46 (.A(sel_R_DATA_TEMPR32[11] ), .B(sel_R_DATA_TEMPR33[11] ), .C(sel_R_DATA_TEMPR34[11] ), .D(sel_R_DATA_TEMPR35[11] ), .Y(OR4_46_Y));
    OR4 OR4_569 (.A(OR4_596_Y), .B(OR4_383_Y), .C(OR4_133_Y), .D(
        OR4_688_Y), .Y(OR4_569_Y));
    OR4 OR4_97 (.A(sel_R_DATA_TEMPR88[12] ), .B(sel_R_DATA_TEMPR89[12] ), .C(sel_R_DATA_TEMPR90[12] ), .D(sel_R_DATA_TEMPR91[12] ), .Y(OR4_97_Y));
    OR4 \OR4_R_DATA[6]  (.A(OR4_323_Y), .B(OR4_977_Y), .C(OR4_51_Y), 
        .D(OR4_243_Y), .Y(R_DATA[6]));
    OR4 OR4_592 (.A(OR4_1036_Y), .B(OR4_534_Y), .C(OR4_1206_Y), .D(
        OR4_678_Y), .Y(OR4_592_Y));
    OR4 OR4_63 (.A(sel_R_DATA_TEMPR52[5] ), .B(sel_R_DATA_TEMPR53[5] ), .C(sel_R_DATA_TEMPR54[5] ), .D(sel_R_DATA_TEMPR55[5] ), .Y(OR4_63_Y));
    OR4 OR4_885 (.A(sel_R_DATA_TEMPR52[20] ), .B(sel_R_DATA_TEMPR53[20] ), 
        .C(sel_R_DATA_TEMPR54[20] ), .D(sel_R_DATA_TEMPR55[20] ), .Y(
        OR4_885_Y));
    OR4 OR4_560 (.A(sel_R_DATA_TEMPR124[10] ), .B(sel_R_DATA_TEMPR125[10] ), 
        .C(sel_R_DATA_TEMPR126[10] ), .D(sel_R_DATA_TEMPR127[10] ), .Y(
        OR4_560_Y));
    OR4 OR4_217 (.A(sel_R_DATA_TEMPR12[26] ), .B(sel_R_DATA_TEMPR13[26] ), 
        .C(sel_R_DATA_TEMPR14[26] ), .D(sel_R_DATA_TEMPR15[26] ), .Y(
        OR4_217_Y));
    OR4 OR4_240 (.A(\SB_CORRECT[28] ), .B(\SB_CORRECT[29] ), .C(
        \SB_CORRECT[30] ), .D(\SB_CORRECT[31] ), .Y(OR4_240_Y));
    OR4 OR4_304 (.A(sel_R_DATA_TEMPR88[15] ), .B(sel_R_DATA_TEMPR89[15] ), 
        .C(sel_R_DATA_TEMPR90[15] ), .D(sel_R_DATA_TEMPR91[15] ), .Y(
        OR4_304_Y));
    OR4 OR4_117 (.A(sel_R_DATA_TEMPR52[27] ), .B(sel_R_DATA_TEMPR53[27] ), 
        .C(sel_R_DATA_TEMPR54[27] ), .D(sel_R_DATA_TEMPR55[27] ), .Y(
        OR4_117_Y));
    OR4 OR4_1203 (.A(OR4_4_Y), .B(OR4_499_Y), .C(OR4_1168_Y), .D(
        OR4_1389_Y), .Y(OR4_1203_Y));
    OR4 OR4_547 (.A(sel_R_DATA_TEMPR104[18] ), .B(sel_R_DATA_TEMPR105[18] ), 
        .C(sel_R_DATA_TEMPR106[18] ), .D(sel_R_DATA_TEMPR107[18] ), .Y(
        OR4_547_Y));
    OR4 OR4_828 (.A(sel_R_DATA_TEMPR20[28] ), .B(sel_R_DATA_TEMPR21[28] ), 
        .C(sel_R_DATA_TEMPR22[28] ), .D(sel_R_DATA_TEMPR23[28] ), .Y(
        OR4_828_Y));
    OR4 OR4_335 (.A(OR4_398_Y), .B(OR4_267_Y), .C(OR4_369_Y), .D(
        OR4_819_Y), .Y(OR4_335_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[3]  (.A(CFG3_19_Y), .B(CFG3_2_Y)
        , .Y(\BLKY2[3] ));
    OR4 OR4_1225 (.A(sel_R_DATA_TEMPR68[5] ), .B(sel_R_DATA_TEMPR69[5] ), .C(sel_R_DATA_TEMPR70[5] ), .D(sel_R_DATA_TEMPR71[5] ), .Y(OR4_1225_Y));
    OR4 \OR4_R_DATA[1]  (.A(OR4_1122_Y), .B(OR4_1299_Y), .C(OR4_912_Y), 
        .D(OR4_724_Y), .Y(R_DATA[1]));
    OR4 OR4_374 (.A(OR4_986_Y), .B(OR4_1227_Y), .C(OR4_1385_Y), .D(
        OR4_705_Y), .Y(OR4_374_Y));
    OR4 OR4_101 (.A(sel_R_DATA_TEMPR64[11] ), .B(sel_R_DATA_TEMPR65[11] ), 
        .C(sel_R_DATA_TEMPR66[11] ), .D(sel_R_DATA_TEMPR67[11] ), .Y(
        OR4_101_Y));
    OR4 OR4_759 (.A(OR4_925_Y), .B(OR4_820_Y), .C(OR4_1289_Y), .D(
        OR4_291_Y), .Y(OR4_759_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[29]  (.A(CFG3_11_Y), .B(
        CFG3_3_Y), .Y(\BLKY2[29] ));
    OR4 OR4_649 (.A(\DB_DETECT[12] ), .B(\DB_DETECT[13] ), .C(
        \DB_DETECT[14] ), .D(\DB_DETECT[15] ), .Y(OR4_649_Y));
    OR4 OR4_594 (.A(sel_R_DATA_TEMPR100[31] ), .B(sel_R_DATA_TEMPR101[31] ), 
        .C(sel_R_DATA_TEMPR102[31] ), .D(sel_R_DATA_TEMPR103[31] ), .Y(
        OR4_594_Y));
    OR4 OR4_171 (.A(sel_R_DATA_TEMPR4[2] ), .B(sel_R_DATA_TEMPR5[2] ), .C(sel_R_DATA_TEMPR6[2] ), .D(sel_R_DATA_TEMPR7[2] ), .Y(OR4_171_Y));
    OR4 OR4_854 (.A(OR4_65_Y), .B(OR4_322_Y), .C(OR4_1251_Y), .D(
        OR4_572_Y), .Y(OR4_854_Y));
    OR4 OR4_1349 (.A(sel_R_DATA_TEMPR120[20] ), .B(sel_R_DATA_TEMPR121[20] ), 
        .C(sel_R_DATA_TEMPR122[20] ), .D(sel_R_DATA_TEMPR123[20] ), .Y(
        OR4_1349_Y));
    OR4 OR4_713 (.A(OR4_1082_Y), .B(OR4_861_Y), .C(OR4_1340_Y), .D(
        OR4_812_Y), .Y(OR4_713_Y));
    OR4 OR4_992 (.A(OR4_1262_Y), .B(OR4_677_Y), .C(OR4_962_Y), .D(
        OR4_286_Y), .Y(OR4_992_Y));
    OR4 OR4_553 (.A(\DB_DETECT[92] ), .B(\DB_DETECT[93] ), .C(
        \DB_DETECT[94] ), .D(\DB_DETECT[95] ), .Y(OR4_553_Y));
    OR4 OR4_1092 (.A(sel_R_DATA_TEMPR108[21] ), .B(sel_R_DATA_TEMPR109[21] ), 
        .C(sel_R_DATA_TEMPR110[21] ), .D(sel_R_DATA_TEMPR111[21] ), .Y(
        OR4_1092_Y));
    OR4 OR4_1040 (.A(sel_R_DATA_TEMPR28[3] ), .B(sel_R_DATA_TEMPR29[3] ), .C(sel_R_DATA_TEMPR30[3] ), .D(sel_R_DATA_TEMPR31[3] ), .Y(OR4_1040_Y));
    OR4 OR4_214 (.A(sel_R_DATA_TEMPR8[1] ), .B(sel_R_DATA_TEMPR9[1] ), .C(sel_R_DATA_TEMPR10[1] ), .D(sel_R_DATA_TEMPR11[1] ), .Y(OR4_214_Y));
    AND4 \AND4SB_CORRECT[45]  (.A(sel_SB_CORRECT_NG[45] ), .B(
        \BLKY2_pipe[11] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[45] ));
    AND4 \AND4SB_CORRECT[46]  (.A(sel_SB_CORRECT_NG[46] ), .B(
        \BLKY2_pipe[11] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[46] ));
    OR4 OR4_246 (.A(sel_R_DATA_TEMPR24[27] ), .B(sel_R_DATA_TEMPR25[27] ), 
        .C(sel_R_DATA_TEMPR26[27] ), .D(sel_R_DATA_TEMPR27[27] ), .Y(
        OR4_246_Y));
    OR4 OR4_221 (.A(OR4_985_Y), .B(OR4_1225_Y), .C(OR4_1384_Y), .D(
        OR4_1185_Y), .Y(OR4_221_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%53%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R53C0 (.A_DOUT({
        nc984, nc985, nc986, nc987, nc988,int_R_DATA_TEMPR53[31] , 
       int_R_DATA_TEMPR53[30] ,int_R_DATA_TEMPR53[29] , 
       int_R_DATA_TEMPR53[28] ,int_R_DATA_TEMPR53[27] , 
       int_R_DATA_TEMPR53[26] ,int_R_DATA_TEMPR53[25] , 
       int_R_DATA_TEMPR53[24] ,int_R_DATA_TEMPR53[23] , 
       int_R_DATA_TEMPR53[22] ,int_R_DATA_TEMPR53[21] , 
       int_R_DATA_TEMPR53[20] ,int_R_DATA_TEMPR53[19] , 
       int_R_DATA_TEMPR53[18] ,int_R_DATA_TEMPR53[17] }), .B_DOUT({nc989, 
        nc990, nc991,int_R_DATA_TEMPR53[16] ,int_R_DATA_TEMPR53[15] , 
       int_R_DATA_TEMPR53[14] ,int_R_DATA_TEMPR53[13] , 
       int_R_DATA_TEMPR53[12] ,int_R_DATA_TEMPR53[11] , 
       int_R_DATA_TEMPR53[10] ,int_R_DATA_TEMPR53[9] ,int_R_DATA_TEMPR53[8] , 
       int_R_DATA_TEMPR53[7] ,int_R_DATA_TEMPR53[6] ,int_R_DATA_TEMPR53[5] , 
       int_R_DATA_TEMPR53[4] ,int_R_DATA_TEMPR53[3] ,int_R_DATA_TEMPR53[2] , 
       int_R_DATA_TEMPR53[1] ,int_R_DATA_TEMPR53[0] }), .DB_DETECT( int_DB_DETECT_NG[53] ), .SB_CORRECT(int_SB_CORRECT_NG[53] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[53] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[13] , \BLKY1[0] , R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[13] , \BLKX1[0] , 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_401 (.A(OR4_638_Y), .B(OR4_506_Y), .C(OR4_600_Y), .D(
        OR4_1201_Y), .Y(OR4_401_Y));
    AND4 \AND4DB_DETECT[99]  (.A(sel_DB_DETECT_NG[99] ), .B(
        \BLKY2_pipe[24] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[99] ));
    OR4 OR4_1109 (.A(sel_R_DATA_TEMPR76[20] ), .B(sel_R_DATA_TEMPR77[20] ), 
        .C(sel_R_DATA_TEMPR78[20] ), .D(sel_R_DATA_TEMPR79[20] ), .Y(
        OR4_1109_Y));
    OR4 OR4_74 (.A(sel_R_DATA_TEMPR64[17] ), .B(sel_R_DATA_TEMPR65[17] ), .C(sel_R_DATA_TEMPR66[17] ), .D(sel_R_DATA_TEMPR67[17] ), .Y(OR4_74_Y));
    OR4 OR4_408 (.A(OR4_53_Y), .B(OR4_708_Y), .C(OR4_1112_Y), .D(
        OR4_1377_Y), .Y(OR4_408_Y));
    OR4 OR4_1283 (.A(sel_R_DATA_TEMPR12[3] ), .B(sel_R_DATA_TEMPR13[3] ), .C(sel_R_DATA_TEMPR14[3] ), .D(sel_R_DATA_TEMPR15[3] ), .Y(OR4_1283_Y));
    OR4 OR4_1259 (.A(sel_R_DATA_TEMPR120[2] ), .B(sel_R_DATA_TEMPR121[2] ), 
        .C(sel_R_DATA_TEMPR122[2] ), .D(sel_R_DATA_TEMPR123[2] ), .Y(
        OR4_1259_Y));
    OR4 OR4_732 (.A(sel_R_DATA_TEMPR56[14] ), .B(sel_R_DATA_TEMPR57[14] ), 
        .C(sel_R_DATA_TEMPR58[14] ), .D(sel_R_DATA_TEMPR59[14] ), .Y(
        OR4_732_Y));
    OR4 OR4_471 (.A(sel_R_DATA_TEMPR72[26] ), .B(sel_R_DATA_TEMPR73[26] ), 
        .C(sel_R_DATA_TEMPR74[26] ), .D(sel_R_DATA_TEMPR75[26] ), .Y(
        OR4_471_Y));
    OR4 OR4_363 (.A(sel_R_DATA_TEMPR16[18] ), .B(sel_R_DATA_TEMPR17[18] ), 
        .C(sel_R_DATA_TEMPR18[18] ), .D(sel_R_DATA_TEMPR19[18] ), .Y(
        OR4_363_Y));
    AND4 \AND4SB_CORRECT[89]  (.A(sel_SB_CORRECT_NG[89] ), .B(
        \BLKY2_pipe[22] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\SB_CORRECT[89] ));
    OR4 OR4_760 (.A(sel_R_DATA_TEMPR88[17] ), .B(sel_R_DATA_TEMPR89[17] ), 
        .C(sel_R_DATA_TEMPR90[17] ), .D(sel_R_DATA_TEMPR91[17] ), .Y(
        OR4_760_Y));
    OR4 OR4_478 (.A(sel_R_DATA_TEMPR12[1] ), .B(sel_R_DATA_TEMPR13[1] ), .C(sel_R_DATA_TEMPR14[1] ), .D(sel_R_DATA_TEMPR15[1] ), .Y(OR4_478_Y));
    OR4 OR4_391 (.A(sel_R_DATA_TEMPR60[2] ), .B(sel_R_DATA_TEMPR61[2] ), .C(sel_R_DATA_TEMPR62[2] ), .D(sel_R_DATA_TEMPR63[2] ), .Y(OR4_391_Y));
    OR4 OR4_936 (.A(OR4_287_Y), .B(OR2_24_Y), .C(sel_R_DATA_TEMPR86[19] ), 
        .D(sel_R_DATA_TEMPR87[19] ), .Y(OR4_936_Y));
    OR4 OR4_644 (.A(sel_R_DATA_TEMPR76[12] ), .B(sel_R_DATA_TEMPR77[12] ), 
        .C(sel_R_DATA_TEMPR78[12] ), .D(sel_R_DATA_TEMPR79[12] ), .Y(
        OR4_644_Y));
    OR4 OR4_61 (.A(sel_R_DATA_TEMPR72[2] ), .B(sel_R_DATA_TEMPR73[2] ), .C(sel_R_DATA_TEMPR74[2] ), .D(sel_R_DATA_TEMPR75[2] ), .Y(OR4_61_Y));
    AND4 \AND4DB_DETECT[69]  (.A(sel_DB_DETECT_NG[69] ), .B(
        \BLKY2_pipe[17] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[0] ), 
        .Y(\DB_DETECT[69] ));
    OR4 OR4_462 (.A(sel_R_DATA_TEMPR88[29] ), .B(sel_R_DATA_TEMPR89[29] ), 
        .C(sel_R_DATA_TEMPR90[29] ), .D(sel_R_DATA_TEMPR91[29] ), .Y(
        OR4_462_Y));
    OR4 OR4_1034 (.A(sel_R_DATA_TEMPR12[24] ), .B(sel_R_DATA_TEMPR13[24] ), 
        .C(sel_R_DATA_TEMPR14[24] ), .D(sel_R_DATA_TEMPR15[24] ), .Y(
        OR4_1034_Y));
    OR4 OR4_635 (.A(sel_R_DATA_TEMPR4[28] ), .B(sel_R_DATA_TEMPR5[28] ), .C(sel_R_DATA_TEMPR6[28] ), .D(sel_R_DATA_TEMPR7[28] ), .Y(OR4_635_Y));
    OR4 OR4_522 (.A(sel_R_DATA_TEMPR44[25] ), .B(sel_R_DATA_TEMPR45[25] ), 
        .C(sel_R_DATA_TEMPR46[25] ), .D(sel_R_DATA_TEMPR47[25] ), .Y(
        OR4_522_Y));
    OR4 OR4_686 (.A(OR4_210_Y), .B(OR4_297_Y), .C(OR4_733_Y), .D(
        OR4_284_Y), .Y(OR4_686_Y));
    AND4 \AND4DB_DETECT[2]  (.A(sel_DB_DETECT_NG[2] ), .B(
        \BLKY2_pipe[0] ), .C(\BLKY0_pipe[0] ), .D(\BLKY1_pipe[1] ), .Y(
        \DB_DETECT[2] ));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%86%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R86C0 (.A_DOUT({
        nc992, nc993, nc994, nc995, nc996,int_R_DATA_TEMPR86[31] , 
       int_R_DATA_TEMPR86[30] ,int_R_DATA_TEMPR86[29] , 
       int_R_DATA_TEMPR86[28] ,int_R_DATA_TEMPR86[27] , 
       int_R_DATA_TEMPR86[26] ,int_R_DATA_TEMPR86[25] , 
       int_R_DATA_TEMPR86[24] ,int_R_DATA_TEMPR86[23] , 
       int_R_DATA_TEMPR86[22] ,int_R_DATA_TEMPR86[21] , 
       int_R_DATA_TEMPR86[20] ,int_R_DATA_TEMPR86[19] , 
       int_R_DATA_TEMPR86[18] ,int_R_DATA_TEMPR86[17] }), .B_DOUT({nc997, 
        nc998, nc999,int_R_DATA_TEMPR86[16] ,int_R_DATA_TEMPR86[15] , 
       int_R_DATA_TEMPR86[14] ,int_R_DATA_TEMPR86[13] , 
       int_R_DATA_TEMPR86[12] ,int_R_DATA_TEMPR86[11] , 
       int_R_DATA_TEMPR86[10] ,int_R_DATA_TEMPR86[9] ,int_R_DATA_TEMPR86[8] , 
       int_R_DATA_TEMPR86[7] ,int_R_DATA_TEMPR86[6] ,int_R_DATA_TEMPR86[5] , 
       int_R_DATA_TEMPR86[4] ,int_R_DATA_TEMPR86[3] ,int_R_DATA_TEMPR86[2] , 
       int_R_DATA_TEMPR86[1] ,int_R_DATA_TEMPR86[0] }), .DB_DETECT( int_DB_DETECT_NG[86] ), .SB_CORRECT(int_SB_CORRECT_NG[86] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[86] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[21] , R_ADDR[10], \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[21] , W_ADDR[10], 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_469 (.A(sel_R_DATA_TEMPR20[31] ), .B(sel_R_DATA_TEMPR21[31] ), 
        .C(sel_R_DATA_TEMPR22[31] ), .D(sel_R_DATA_TEMPR23[31] ), .Y(
        OR4_469_Y));
    OR2 OR2_5 (.A(sel_R_DATA_TEMPR84[3] ), .B(sel_R_DATA_TEMPR85[3] ), .Y(
        OR2_5_Y));
    OR4 OR4_315 (.A(OR4_392_Y), .B(OR4_1306_Y), .C(OR4_674_Y), .D(
        OR4_612_Y), .Y(OR4_315_Y));
    OR4 OR4_1333 (.A(sel_R_DATA_TEMPR92[29] ), .B(sel_R_DATA_TEMPR93[29] ), 
        .C(sel_R_DATA_TEMPR94[29] ), .D(sel_R_DATA_TEMPR95[29] ), .Y(
        OR4_1333_Y));
    OR4 OR4_490 (.A(sel_R_DATA_TEMPR0[16] ), .B(sel_R_DATA_TEMPR1[16] ), .C(sel_R_DATA_TEMPR2[16] ), .D(sel_R_DATA_TEMPR3[16] ), .Y(OR4_490_Y));
    OR4 OR4_40 (.A(sel_R_DATA_TEMPR124[23] ), .B(sel_R_DATA_TEMPR125[23] ), 
        .C(sel_R_DATA_TEMPR126[23] ), .D(sel_R_DATA_TEMPR127[23] ), .Y(
        OR4_40_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%11%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R11C0 (.A_DOUT({
        nc1000, nc1001, nc1002, nc1003, nc1004,int_R_DATA_TEMPR11[31] , 
       int_R_DATA_TEMPR11[30] ,int_R_DATA_TEMPR11[29] , 
       int_R_DATA_TEMPR11[28] ,int_R_DATA_TEMPR11[27] , 
       int_R_DATA_TEMPR11[26] ,int_R_DATA_TEMPR11[25] , 
       int_R_DATA_TEMPR11[24] ,int_R_DATA_TEMPR11[23] , 
       int_R_DATA_TEMPR11[22] ,int_R_DATA_TEMPR11[21] , 
       int_R_DATA_TEMPR11[20] ,int_R_DATA_TEMPR11[19] , 
       int_R_DATA_TEMPR11[18] ,int_R_DATA_TEMPR11[17] }), .B_DOUT({nc1005, 
        nc1006, nc1007,int_R_DATA_TEMPR11[16] ,int_R_DATA_TEMPR11[15] , 
       int_R_DATA_TEMPR11[14] ,int_R_DATA_TEMPR11[13] , 
       int_R_DATA_TEMPR11[12] ,int_R_DATA_TEMPR11[11] , 
       int_R_DATA_TEMPR11[10] ,int_R_DATA_TEMPR11[9] ,int_R_DATA_TEMPR11[8] , 
       int_R_DATA_TEMPR11[7] ,int_R_DATA_TEMPR11[6] ,int_R_DATA_TEMPR11[5] , 
       int_R_DATA_TEMPR11[4] ,int_R_DATA_TEMPR11[3] ,int_R_DATA_TEMPR11[2] , 
       int_R_DATA_TEMPR11[1] ,int_R_DATA_TEMPR11[0] }), .DB_DETECT( int_DB_DETECT_NG[11] ), .SB_CORRECT(int_SB_CORRECT_NG[11] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[11] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[2] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[2] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_509 (.A(sel_R_DATA_TEMPR92[22] ), .B(sel_R_DATA_TEMPR93[22] ), 
        .C(sel_R_DATA_TEMPR94[22] ), .D(sel_R_DATA_TEMPR95[22] ), .Y(
        OR4_509_Y));
    OR4 OR4_166 (.A(sel_R_DATA_TEMPR120[4] ), .B(sel_R_DATA_TEMPR121[4] ), 
        .C(sel_R_DATA_TEMPR122[4] ), .D(sel_R_DATA_TEMPR123[4] ), .Y(
        OR4_166_Y));
    OR4 OR4_1189 (.A(sel_R_DATA_TEMPR32[2] ), .B(sel_R_DATA_TEMPR33[2] ), .C(sel_R_DATA_TEMPR34[2] ), .D(sel_R_DATA_TEMPR35[2] ), .Y(OR4_1189_Y));
    CFG2 #( .INIT(4'h8) )  \CFG2_BLKY2[26]  (.A(CFG3_0_Y), .B(CFG3_3_Y)
        , .Y(\BLKY2[26] ));
    OR4 OR4_500 (.A(sel_R_DATA_TEMPR12[5] ), .B(sel_R_DATA_TEMPR13[5] ), .C(sel_R_DATA_TEMPR14[5] ), .D(sel_R_DATA_TEMPR15[5] ), .Y(OR4_500_Y));
    AND4 \AND4SB_CORRECT[115]  (.A(sel_SB_CORRECT_NG[115] ), .B(
        \BLKY2_pipe[28] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\SB_CORRECT[115] ));
    OR4 OR4_47 (.A(sel_R_DATA_TEMPR24[5] ), .B(sel_R_DATA_TEMPR25[5] ), .C(sel_R_DATA_TEMPR26[5] ), .D(sel_R_DATA_TEMPR27[5] ), .Y(OR4_47_Y));
    OR4 OR4_1106 (.A(sel_R_DATA_TEMPR64[23] ), .B(sel_R_DATA_TEMPR65[23] ), 
        .C(sel_R_DATA_TEMPR66[23] ), .D(sel_R_DATA_TEMPR67[23] ), .Y(
        OR4_1106_Y));
    OR4 OR4_579 (.A(sel_R_DATA_TEMPR20[19] ), .B(sel_R_DATA_TEMPR21[19] ), 
        .C(sel_R_DATA_TEMPR22[19] ), .D(sel_R_DATA_TEMPR23[19] ), .Y(
        OR4_579_Y));
    OR4 OR4_1113 (.A(sel_R_DATA_TEMPR8[12] ), .B(sel_R_DATA_TEMPR9[12] ), .C(sel_R_DATA_TEMPR10[12] ), .D(sel_R_DATA_TEMPR11[12] ), .Y(OR4_1113_Y)
        );
    OR4 OR4_570 (.A(sel_R_DATA_TEMPR48[13] ), .B(sel_R_DATA_TEMPR49[13] ), 
        .C(sel_R_DATA_TEMPR50[13] ), .D(sel_R_DATA_TEMPR51[13] ), .Y(
        OR4_570_Y));
    OR4 OR4_1375 (.A(sel_R_DATA_TEMPR40[5] ), .B(sel_R_DATA_TEMPR41[5] ), .C(sel_R_DATA_TEMPR42[5] ), .D(sel_R_DATA_TEMPR43[5] ), .Y(OR4_1375_Y));
    OR4 OR4_524 (.A(sel_R_DATA_TEMPR80[17] ), .B(sel_R_DATA_TEMPR81[17] ), 
        .C(sel_R_DATA_TEMPR82[17] ), .D(sel_R_DATA_TEMPR83[17] ), .Y(
        OR4_524_Y));
    OR4 OR4_1201 (.A(sel_R_DATA_TEMPR76[18] ), .B(sel_R_DATA_TEMPR77[18] ), 
        .C(sel_R_DATA_TEMPR78[18] ), .D(sel_R_DATA_TEMPR79[18] ), .Y(
        OR4_1201_Y));
    OR4 OR4_1108 (.A(sel_R_DATA_TEMPR96[21] ), .B(sel_R_DATA_TEMPR97[21] ), 
        .C(sel_R_DATA_TEMPR98[21] ), .D(sel_R_DATA_TEMPR99[21] ), .Y(
        OR4_1108_Y));
    OR4 \OR4_R_DATA[28]  (.A(OR4_1214_Y), .B(OR4_1013_Y), .C(OR4_385_Y)
        , .D(OR4_569_Y), .Y(R_DATA[28]));
    OR4 OR4_922 (.A(OR4_1060_Y), .B(OR4_1290_Y), .C(OR4_61_Y), .D(
        OR4_1074_Y), .Y(OR4_922_Y));
    OR4 OR4_368 (.A(OR4_111_Y), .B(OR4_410_Y), .C(OR4_851_Y), .D(
        OR4_350_Y), .Y(OR4_368_Y));
    OR4 OR4_712 (.A(sel_R_DATA_TEMPR4[12] ), .B(sel_R_DATA_TEMPR5[12] ), .C(sel_R_DATA_TEMPR6[12] ), .D(sel_R_DATA_TEMPR7[12] ), .Y(OR4_712_Y));
    AND4 \AND4DB_DETECT[107]  (.A(sel_DB_DETECT_NG[107] ), .B(
        \BLKY2_pipe[26] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[107] ));
    OR4 OR4_630 (.A(sel_R_DATA_TEMPR52[23] ), .B(sel_R_DATA_TEMPR53[23] ), 
        .C(sel_R_DATA_TEMPR54[23] ), .D(sel_R_DATA_TEMPR55[23] ), .Y(
        OR4_630_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%20%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R20C0 (.A_DOUT({
        nc1008, nc1009, nc1010, nc1011, nc1012,int_R_DATA_TEMPR20[31] , 
       int_R_DATA_TEMPR20[30] ,int_R_DATA_TEMPR20[29] , 
       int_R_DATA_TEMPR20[28] ,int_R_DATA_TEMPR20[27] , 
       int_R_DATA_TEMPR20[26] ,int_R_DATA_TEMPR20[25] , 
       int_R_DATA_TEMPR20[24] ,int_R_DATA_TEMPR20[23] , 
       int_R_DATA_TEMPR20[22] ,int_R_DATA_TEMPR20[21] , 
       int_R_DATA_TEMPR20[20] ,int_R_DATA_TEMPR20[19] , 
       int_R_DATA_TEMPR20[18] ,int_R_DATA_TEMPR20[17] }), .B_DOUT({nc1013, 
        nc1014, nc1015,int_R_DATA_TEMPR20[16] ,int_R_DATA_TEMPR20[15] , 
       int_R_DATA_TEMPR20[14] ,int_R_DATA_TEMPR20[13] , 
       int_R_DATA_TEMPR20[12] ,int_R_DATA_TEMPR20[11] , 
       int_R_DATA_TEMPR20[10] ,int_R_DATA_TEMPR20[9] ,int_R_DATA_TEMPR20[8] , 
       int_R_DATA_TEMPR20[7] ,int_R_DATA_TEMPR20[6] ,int_R_DATA_TEMPR20[5] , 
       int_R_DATA_TEMPR20[4] ,int_R_DATA_TEMPR20[3] ,int_R_DATA_TEMPR20[2] , 
       int_R_DATA_TEMPR20[1] ,int_R_DATA_TEMPR20[0] }), .DB_DETECT( int_DB_DETECT_NG[20] ), .SB_CORRECT(int_SB_CORRECT_NG[20] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[20] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[5] , \BLKY1[0] , \BLKY0[0] }), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[5] , \BLKX1[0] , 
        \BLKX0[0] }), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    AND4 \AND4DB_DETECT[43]  (.A(sel_DB_DETECT_NG[43] ), .B(
        \BLKY2_pipe[10] ), .C(\BLKY0_pipe[1] ), .D(\BLKY1_pipe[1] ), 
        .Y(\DB_DETECT[43] ));
    OR4 OR4_916 (.A(sel_R_DATA_TEMPR44[6] ), .B(sel_R_DATA_TEMPR45[6] ), .C(sel_R_DATA_TEMPR46[6] ), .D(sel_R_DATA_TEMPR47[6] ), .Y(OR4_916_Y));
    OR4 OR4_98 (.A(sel_R_DATA_TEMPR32[6] ), .B(sel_R_DATA_TEMPR33[6] ), .C(sel_R_DATA_TEMPR34[6] ), .D(sel_R_DATA_TEMPR35[6] ), .Y(OR4_98_Y));
    RAM1K20 #( .RAMINDEX("PF_TPSRAM_MAX_0%65536-65536%32-32%POWER%119%0%TWO-PORT%ECC_EN-2")
         )  miv_rv32_ram_singleport_lp_ecc_R119C0 (.A_DOUT({
        nc1016, nc1017, nc1018, nc1019, nc1020,int_R_DATA_TEMPR119[31] , 
       int_R_DATA_TEMPR119[30] ,int_R_DATA_TEMPR119[29] , 
       int_R_DATA_TEMPR119[28] ,int_R_DATA_TEMPR119[27] , 
       int_R_DATA_TEMPR119[26] ,int_R_DATA_TEMPR119[25] , 
       int_R_DATA_TEMPR119[24] ,int_R_DATA_TEMPR119[23] , 
       int_R_DATA_TEMPR119[22] ,int_R_DATA_TEMPR119[21] , 
       int_R_DATA_TEMPR119[20] ,int_R_DATA_TEMPR119[19] , 
       int_R_DATA_TEMPR119[18] ,int_R_DATA_TEMPR119[17] }), .B_DOUT({
        nc1021, nc1022, nc1023,int_R_DATA_TEMPR119[16] , 
       int_R_DATA_TEMPR119[15] ,int_R_DATA_TEMPR119[14] , 
       int_R_DATA_TEMPR119[13] ,int_R_DATA_TEMPR119[12] , 
       int_R_DATA_TEMPR119[11] ,int_R_DATA_TEMPR119[10] , 
       int_R_DATA_TEMPR119[9] ,int_R_DATA_TEMPR119[8] , 
       int_R_DATA_TEMPR119[7] ,int_R_DATA_TEMPR119[6] , 
       int_R_DATA_TEMPR119[5] ,int_R_DATA_TEMPR119[4] , 
       int_R_DATA_TEMPR119[3] ,int_R_DATA_TEMPR119[2] , 
       int_R_DATA_TEMPR119[1] ,int_R_DATA_TEMPR119[0] }), .DB_DETECT( int_DB_DETECT_NG[119] ), .SB_CORRECT(int_SB_CORRECT_NG[119] ), 
        .ACCESS_BUSY(\ACCESS_BUSY[119] ), .A_ADDR({R_ADDR[8], 
        R_ADDR[7], R_ADDR[6], R_ADDR[5], R_ADDR[4], R_ADDR[3], 
        R_ADDR[2], R_ADDR[1], R_ADDR[0], GND, GND, GND, GND, GND}), 
        .A_BLK_EN({\BLKY2[29] , R_ADDR[10], R_ADDR[9]}), .A_CLK(CLK), 
        .A_DIN({GND, GND, GND, GND, GND, W_DATA[31], W_DATA[30], 
        W_DATA[29], W_DATA[28], W_DATA[27], W_DATA[26], W_DATA[25], 
        W_DATA[24], W_DATA[23], W_DATA[22], W_DATA[21], W_DATA[20], 
        W_DATA[19], W_DATA[18], W_DATA[17]}), .A_REN(VCC), .A_WEN({VCC, 
        VCC}), .A_DOUT_EN(VCC), .A_DOUT_ARST_N(VCC), .A_DOUT_SRST_N(
        VCC), .B_ADDR({W_ADDR[8], W_ADDR[7], W_ADDR[6], W_ADDR[5], 
        W_ADDR[4], W_ADDR[3], W_ADDR[2], W_ADDR[1], W_ADDR[0], GND, 
        GND, GND, GND, GND}), .B_BLK_EN({\BLKX2[29] , W_ADDR[10], 
        W_ADDR[9]}), .B_CLK(CLK), .B_DIN({GND, GND, GND, W_DATA[16], 
        W_DATA[15], W_DATA[14], W_DATA[13], W_DATA[12], W_DATA[11], 
        W_DATA[10], W_DATA[9], W_DATA[8], W_DATA[7], W_DATA[6], 
        W_DATA[5], W_DATA[4], W_DATA[3], W_DATA[2], W_DATA[1], 
        W_DATA[0]}), .B_REN(VCC), .B_WEN({VCC, VCC}), .B_DOUT_EN(VCC), 
        .B_DOUT_ARST_N(VCC), .B_DOUT_SRST_N(VCC), .ECC_EN(VCC), 
        .BUSY_FB(GND), .A_WIDTH({VCC, GND, VCC}), .A_WMODE({GND, GND}), 
        .A_BYPASS(VCC), .B_WIDTH({VCC, GND, VCC}), .B_WMODE({GND, GND})
        , .B_BYPASS(VCC), .ECC_BYPASS(VCC));
    OR4 OR4_1024 (.A(sel_R_DATA_TEMPR48[27] ), .B(sel_R_DATA_TEMPR49[27] ), 
        .C(sel_R_DATA_TEMPR50[27] ), .D(sel_R_DATA_TEMPR51[27] ), .Y(
        OR4_1024_Y));
    OR4 OR4_321 (.A(OR4_1062_Y), .B(OR4_433_Y), .C(OR4_402_Y), .D(
        OR4_1059_Y), .Y(OR4_321_Y));
    OR4 OR4_1186 (.A(sel_R_DATA_TEMPR88[8] ), .B(sel_R_DATA_TEMPR89[8] ), .C(sel_R_DATA_TEMPR90[8] ), .D(sel_R_DATA_TEMPR91[8] ), .Y(OR4_1186_Y));
    OR4 OR4_615 (.A(sel_R_DATA_TEMPR36[14] ), .B(sel_R_DATA_TEMPR37[14] ), 
        .C(sel_R_DATA_TEMPR38[14] ), .D(sel_R_DATA_TEMPR39[14] ), .Y(
        OR4_615_Y));
    OR4 OR4_337 (.A(sel_R_DATA_TEMPR4[24] ), .B(sel_R_DATA_TEMPR5[24] ), .C(sel_R_DATA_TEMPR6[24] ), .D(sel_R_DATA_TEMPR7[24] ), .Y(OR4_337_Y));
    OR4 OR4_130 (.A(sel_R_DATA_TEMPR120[24] ), .B(sel_R_DATA_TEMPR121[24] ), 
        .C(sel_R_DATA_TEMPR122[24] ), .D(sel_R_DATA_TEMPR123[24] ), .Y(
        OR4_130_Y));
    OR2 OR2_25 (.A(sel_R_DATA_TEMPR84[22] ), .B(sel_R_DATA_TEMPR85[22] ), .Y(
        OR2_25_Y));
    OR4 OR4_1323 (.A(sel_R_DATA_TEMPR100[2] ), .B(sel_R_DATA_TEMPR101[2] ), 
        .C(sel_R_DATA_TEMPR102[2] ), .D(sel_R_DATA_TEMPR103[2] ), .Y(
        OR4_1323_Y));
    OR4 OR4_1036 (.A(\DB_DETECT[96] ), .B(\DB_DETECT[97] ), .C(
        \DB_DETECT[98] ), .D(\DB_DETECT[99] ), .Y(OR4_1036_Y));
    OR4 OR4_1281 (.A(sel_R_DATA_TEMPR112[10] ), .B(sel_R_DATA_TEMPR113[10] ), 
        .C(sel_R_DATA_TEMPR114[10] ), .D(sel_R_DATA_TEMPR115[10] ), .Y(
        OR4_1281_Y));
    OR4 OR4_169 (.A(sel_R_DATA_TEMPR80[9] ), .B(sel_R_DATA_TEMPR81[9] ), .C(sel_R_DATA_TEMPR82[9] ), .D(sel_R_DATA_TEMPR83[9] ), .Y(OR4_169_Y));
    OR4 OR4_303 (.A(OR4_199_Y), .B(OR4_1382_Y), .C(OR4_180_Y), .D(
        OR4_1161_Y), .Y(OR4_303_Y));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
